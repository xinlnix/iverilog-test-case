module mux4_1();
    input in0, in1, in2, in3;
    input [1:0] sel;
    integer i;

    reg [7:0] out1;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1 = in0;
    end

    reg [7:0] out2;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2 = in0;
    end

    reg [7:0] out3;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3 = in0;
    end

    reg [7:0] out4;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4 = in0;
    end

    reg [7:0] out5;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5 = in0;
    end

    reg [7:0] out6;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6 = in0;
    end

    reg [7:0] out7;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7 = in0;
    end

    reg [7:0] out8;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8 = in0;
    end

    reg [7:0] out9;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9 = in0;
    end

    reg [7:0] out10;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out10 = in0;
    end

    reg [7:0] out11;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out11 = in0;
    end

    reg [7:0] out12;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out12 = in0;
    end

    reg [7:0] out13;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out13 = in0;
    end

    reg [7:0] out14;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out14 = in0;
    end

    reg [7:0] out15;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out15 = in0;
    end

    reg [7:0] out16;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out16 = in0;
    end

    reg [7:0] out17;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out17 = in0;
    end

    reg [7:0] out18;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out18 = in0;
    end

    reg [7:0] out19;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out19 = in0;
    end

    reg [7:0] out20;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out20 = in0;
    end

    reg [7:0] out21;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out21 = in0;
    end

    reg [7:0] out22;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out22 = in0;
    end

    reg [7:0] out23;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out23 = in0;
    end

    reg [7:0] out24;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out24 = in0;
    end

    reg [7:0] out25;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out25 = in0;
    end

    reg [7:0] out26;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out26 = in0;
    end

    reg [7:0] out27;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out27 = in0;
    end

    reg [7:0] out28;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out28 = in0;
    end

    reg [7:0] out29;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out29 = in0;
    end

    reg [7:0] out30;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out30 = in0;
    end

    reg [7:0] out31;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out31 = in0;
    end

    reg [7:0] out32;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out32 = in0;
    end

    reg [7:0] out33;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out33 = in0;
    end

    reg [7:0] out34;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out34 = in0;
    end

    reg [7:0] out35;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out35 = in0;
    end

    reg [7:0] out36;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out36 = in0;
    end

    reg [7:0] out37;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out37 = in0;
    end

    reg [7:0] out38;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out38 = in0;
    end

    reg [7:0] out39;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out39 = in0;
    end

    reg [7:0] out40;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out40 = in0;
    end

    reg [7:0] out41;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out41 = in0;
    end

    reg [7:0] out42;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out42 = in0;
    end

    reg [7:0] out43;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out43 = in0;
    end

    reg [7:0] out44;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out44 = in0;
    end

    reg [7:0] out45;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out45 = in0;
    end

    reg [7:0] out46;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out46 = in0;
    end

    reg [7:0] out47;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out47 = in0;
    end

    reg [7:0] out48;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out48 = in0;
    end

    reg [7:0] out49;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out49 = in0;
    end

    reg [7:0] out50;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out50 = in0;
    end

    reg [7:0] out51;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out51 = in0;
    end

    reg [7:0] out52;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out52 = in0;
    end

    reg [7:0] out53;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out53 = in0;
    end

    reg [7:0] out54;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out54 = in0;
    end

    reg [7:0] out55;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out55 = in0;
    end

    reg [7:0] out56;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out56 = in0;
    end

    reg [7:0] out57;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out57 = in0;
    end

    reg [7:0] out58;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out58 = in0;
    end

    reg [7:0] out59;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out59 = in0;
    end

    reg [7:0] out60;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out60 = in0;
    end

    reg [7:0] out61;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out61 = in0;
    end

    reg [7:0] out62;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out62 = in0;
    end

    reg [7:0] out63;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out63 = in0;
    end

    reg [7:0] out64;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out64 = in0;
    end

    reg [7:0] out65;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out65 = in0;
    end

    reg [7:0] out66;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out66 = in0;
    end

    reg [7:0] out67;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out67 = in0;
    end

    reg [7:0] out68;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out68 = in0;
    end

    reg [7:0] out69;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out69 = in0;
    end

    reg [7:0] out70;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out70 = in0;
    end

    reg [7:0] out71;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out71 = in0;
    end

    reg [7:0] out72;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out72 = in0;
    end

    reg [7:0] out73;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out73 = in0;
    end

    reg [7:0] out74;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out74 = in0;
    end

    reg [7:0] out75;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out75 = in0;
    end

    reg [7:0] out76;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out76 = in0;
    end

    reg [7:0] out77;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out77 = in0;
    end

    reg [7:0] out78;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out78 = in0;
    end

    reg [7:0] out79;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out79 = in0;
    end

    reg [7:0] out80;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out80 = in0;
    end

    reg [7:0] out81;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out81 = in0;
    end

    reg [7:0] out82;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out82 = in0;
    end

    reg [7:0] out83;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out83 = in0;
    end

    reg [7:0] out84;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out84 = in0;
    end

    reg [7:0] out85;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out85 = in0;
    end

    reg [7:0] out86;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out86 = in0;
    end

    reg [7:0] out87;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out87 = in0;
    end

    reg [7:0] out88;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out88 = in0;
    end

    reg [7:0] out89;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out89 = in0;
    end

    reg [7:0] out90;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out90 = in0;
    end

    reg [7:0] out91;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out91 = in0;
    end

    reg [7:0] out92;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out92 = in0;
    end

    reg [7:0] out93;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out93 = in0;
    end

    reg [7:0] out94;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out94 = in0;
    end

    reg [7:0] out95;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out95 = in0;
    end

    reg [7:0] out96;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out96 = in0;
    end

    reg [7:0] out97;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out97 = in0;
    end

    reg [7:0] out98;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out98 = in0;
    end

    reg [7:0] out99;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out99 = in0;
    end

    reg [7:0] out100;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out100 = in0;
    end

    reg [7:0] out101;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out101 = in0;
    end

    reg [7:0] out102;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out102 = in0;
    end

    reg [7:0] out103;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out103 = in0;
    end

    reg [7:0] out104;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out104 = in0;
    end

    reg [7:0] out105;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out105 = in0;
    end

    reg [7:0] out106;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out106 = in0;
    end

    reg [7:0] out107;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out107 = in0;
    end

    reg [7:0] out108;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out108 = in0;
    end

    reg [7:0] out109;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out109 = in0;
    end

    reg [7:0] out110;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out110 = in0;
    end

    reg [7:0] out111;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out111 = in0;
    end

    reg [7:0] out112;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out112 = in0;
    end

    reg [7:0] out113;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out113 = in0;
    end

    reg [7:0] out114;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out114 = in0;
    end

    reg [7:0] out115;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out115 = in0;
    end

    reg [7:0] out116;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out116 = in0;
    end

    reg [7:0] out117;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out117 = in0;
    end

    reg [7:0] out118;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out118 = in0;
    end

    reg [7:0] out119;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out119 = in0;
    end

    reg [7:0] out120;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out120 = in0;
    end

    reg [7:0] out121;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out121 = in0;
    end

    reg [7:0] out122;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out122 = in0;
    end

    reg [7:0] out123;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out123 = in0;
    end

    reg [7:0] out124;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out124 = in0;
    end

    reg [7:0] out125;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out125 = in0;
    end

    reg [7:0] out126;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out126 = in0;
    end

    reg [7:0] out127;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out127 = in0;
    end

    reg [7:0] out128;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out128 = in0;
    end

    reg [7:0] out129;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out129 = in0;
    end

    reg [7:0] out130;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out130 = in0;
    end

    reg [7:0] out131;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out131 = in0;
    end

    reg [7:0] out132;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out132 = in0;
    end

    reg [7:0] out133;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out133 = in0;
    end

    reg [7:0] out134;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out134 = in0;
    end

    reg [7:0] out135;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out135 = in0;
    end

    reg [7:0] out136;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out136 = in0;
    end

    reg [7:0] out137;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out137 = in0;
    end

    reg [7:0] out138;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out138 = in0;
    end

    reg [7:0] out139;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out139 = in0;
    end

    reg [7:0] out140;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out140 = in0;
    end

    reg [7:0] out141;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out141 = in0;
    end

    reg [7:0] out142;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out142 = in0;
    end

    reg [7:0] out143;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out143 = in0;
    end

    reg [7:0] out144;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out144 = in0;
    end

    reg [7:0] out145;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out145 = in0;
    end

    reg [7:0] out146;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out146 = in0;
    end

    reg [7:0] out147;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out147 = in0;
    end

    reg [7:0] out148;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out148 = in0;
    end

    reg [7:0] out149;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out149 = in0;
    end

    reg [7:0] out150;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out150 = in0;
    end

    reg [7:0] out151;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out151 = in0;
    end

    reg [7:0] out152;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out152 = in0;
    end

    reg [7:0] out153;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out153 = in0;
    end

    reg [7:0] out154;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out154 = in0;
    end

    reg [7:0] out155;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out155 = in0;
    end

    reg [7:0] out156;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out156 = in0;
    end

    reg [7:0] out157;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out157 = in0;
    end

    reg [7:0] out158;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out158 = in0;
    end

    reg [7:0] out159;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out159 = in0;
    end

    reg [7:0] out160;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out160 = in0;
    end

    reg [7:0] out161;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out161 = in0;
    end

    reg [7:0] out162;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out162 = in0;
    end

    reg [7:0] out163;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out163 = in0;
    end

    reg [7:0] out164;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out164 = in0;
    end

    reg [7:0] out165;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out165 = in0;
    end

    reg [7:0] out166;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out166 = in0;
    end

    reg [7:0] out167;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out167 = in0;
    end

    reg [7:0] out168;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out168 = in0;
    end

    reg [7:0] out169;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out169 = in0;
    end

    reg [7:0] out170;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out170 = in0;
    end

    reg [7:0] out171;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out171 = in0;
    end

    reg [7:0] out172;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out172 = in0;
    end

    reg [7:0] out173;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out173 = in0;
    end

    reg [7:0] out174;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out174 = in0;
    end

    reg [7:0] out175;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out175 = in0;
    end

    reg [7:0] out176;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out176 = in0;
    end

    reg [7:0] out177;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out177 = in0;
    end

    reg [7:0] out178;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out178 = in0;
    end

    reg [7:0] out179;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out179 = in0;
    end

    reg [7:0] out180;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out180 = in0;
    end

    reg [7:0] out181;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out181 = in0;
    end

    reg [7:0] out182;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out182 = in0;
    end

    reg [7:0] out183;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out183 = in0;
    end

    reg [7:0] out184;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out184 = in0;
    end

    reg [7:0] out185;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out185 = in0;
    end

    reg [7:0] out186;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out186 = in0;
    end

    reg [7:0] out187;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out187 = in0;
    end

    reg [7:0] out188;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out188 = in0;
    end

    reg [7:0] out189;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out189 = in0;
    end

    reg [7:0] out190;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out190 = in0;
    end

    reg [7:0] out191;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out191 = in0;
    end

    reg [7:0] out192;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out192 = in0;
    end

    reg [7:0] out193;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out193 = in0;
    end

    reg [7:0] out194;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out194 = in0;
    end

    reg [7:0] out195;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out195 = in0;
    end

    reg [7:0] out196;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out196 = in0;
    end

    reg [7:0] out197;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out197 = in0;
    end

    reg [7:0] out198;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out198 = in0;
    end

    reg [7:0] out199;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out199 = in0;
    end

    reg [7:0] out200;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out200 = in0;
    end

    reg [7:0] out201;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out201 = in0;
    end

    reg [7:0] out202;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out202 = in0;
    end

    reg [7:0] out203;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out203 = in0;
    end

    reg [7:0] out204;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out204 = in0;
    end

    reg [7:0] out205;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out205 = in0;
    end

    reg [7:0] out206;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out206 = in0;
    end

    reg [7:0] out207;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out207 = in0;
    end

    reg [7:0] out208;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out208 = in0;
    end

    reg [7:0] out209;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out209 = in0;
    end

    reg [7:0] out210;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out210 = in0;
    end

    reg [7:0] out211;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out211 = in0;
    end

    reg [7:0] out212;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out212 = in0;
    end

    reg [7:0] out213;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out213 = in0;
    end

    reg [7:0] out214;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out214 = in0;
    end

    reg [7:0] out215;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out215 = in0;
    end

    reg [7:0] out216;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out216 = in0;
    end

    reg [7:0] out217;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out217 = in0;
    end

    reg [7:0] out218;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out218 = in0;
    end

    reg [7:0] out219;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out219 = in0;
    end

    reg [7:0] out220;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out220 = in0;
    end

    reg [7:0] out221;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out221 = in0;
    end

    reg [7:0] out222;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out222 = in0;
    end

    reg [7:0] out223;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out223 = in0;
    end

    reg [7:0] out224;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out224 = in0;
    end

    reg [7:0] out225;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out225 = in0;
    end

    reg [7:0] out226;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out226 = in0;
    end

    reg [7:0] out227;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out227 = in0;
    end

    reg [7:0] out228;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out228 = in0;
    end

    reg [7:0] out229;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out229 = in0;
    end

    reg [7:0] out230;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out230 = in0;
    end

    reg [7:0] out231;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out231 = in0;
    end

    reg [7:0] out232;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out232 = in0;
    end

    reg [7:0] out233;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out233 = in0;
    end

    reg [7:0] out234;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out234 = in0;
    end

    reg [7:0] out235;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out235 = in0;
    end

    reg [7:0] out236;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out236 = in0;
    end

    reg [7:0] out237;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out237 = in0;
    end

    reg [7:0] out238;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out238 = in0;
    end

    reg [7:0] out239;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out239 = in0;
    end

    reg [7:0] out240;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out240 = in0;
    end

    reg [7:0] out241;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out241 = in0;
    end

    reg [7:0] out242;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out242 = in0;
    end

    reg [7:0] out243;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out243 = in0;
    end

    reg [7:0] out244;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out244 = in0;
    end

    reg [7:0] out245;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out245 = in0;
    end

    reg [7:0] out246;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out246 = in0;
    end

    reg [7:0] out247;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out247 = in0;
    end

    reg [7:0] out248;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out248 = in0;
    end

    reg [7:0] out249;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out249 = in0;
    end

    reg [7:0] out250;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out250 = in0;
    end

    reg [7:0] out251;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out251 = in0;
    end

    reg [7:0] out252;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out252 = in0;
    end

    reg [7:0] out253;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out253 = in0;
    end

    reg [7:0] out254;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out254 = in0;
    end

    reg [7:0] out255;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out255 = in0;
    end

    reg [7:0] out256;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out256 = in0;
    end

    reg [7:0] out257;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out257 = in0;
    end

    reg [7:0] out258;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out258 = in0;
    end

    reg [7:0] out259;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out259 = in0;
    end

    reg [7:0] out260;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out260 = in0;
    end

    reg [7:0] out261;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out261 = in0;
    end

    reg [7:0] out262;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out262 = in0;
    end

    reg [7:0] out263;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out263 = in0;
    end

    reg [7:0] out264;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out264 = in0;
    end

    reg [7:0] out265;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out265 = in0;
    end

    reg [7:0] out266;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out266 = in0;
    end

    reg [7:0] out267;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out267 = in0;
    end

    reg [7:0] out268;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out268 = in0;
    end

    reg [7:0] out269;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out269 = in0;
    end

    reg [7:0] out270;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out270 = in0;
    end

    reg [7:0] out271;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out271 = in0;
    end

    reg [7:0] out272;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out272 = in0;
    end

    reg [7:0] out273;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out273 = in0;
    end

    reg [7:0] out274;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out274 = in0;
    end

    reg [7:0] out275;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out275 = in0;
    end

    reg [7:0] out276;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out276 = in0;
    end

    reg [7:0] out277;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out277 = in0;
    end

    reg [7:0] out278;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out278 = in0;
    end

    reg [7:0] out279;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out279 = in0;
    end

    reg [7:0] out280;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out280 = in0;
    end

    reg [7:0] out281;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out281 = in0;
    end

    reg [7:0] out282;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out282 = in0;
    end

    reg [7:0] out283;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out283 = in0;
    end

    reg [7:0] out284;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out284 = in0;
    end

    reg [7:0] out285;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out285 = in0;
    end

    reg [7:0] out286;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out286 = in0;
    end

    reg [7:0] out287;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out287 = in0;
    end

    reg [7:0] out288;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out288 = in0;
    end

    reg [7:0] out289;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out289 = in0;
    end

    reg [7:0] out290;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out290 = in0;
    end

    reg [7:0] out291;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out291 = in0;
    end

    reg [7:0] out292;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out292 = in0;
    end

    reg [7:0] out293;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out293 = in0;
    end

    reg [7:0] out294;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out294 = in0;
    end

    reg [7:0] out295;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out295 = in0;
    end

    reg [7:0] out296;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out296 = in0;
    end

    reg [7:0] out297;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out297 = in0;
    end

    reg [7:0] out298;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out298 = in0;
    end

    reg [7:0] out299;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out299 = in0;
    end

    reg [7:0] out300;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out300 = in0;
    end

    reg [7:0] out301;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out301 = in0;
    end

    reg [7:0] out302;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out302 = in0;
    end

    reg [7:0] out303;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out303 = in0;
    end

    reg [7:0] out304;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out304 = in0;
    end

    reg [7:0] out305;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out305 = in0;
    end

    reg [7:0] out306;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out306 = in0;
    end

    reg [7:0] out307;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out307 = in0;
    end

    reg [7:0] out308;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out308 = in0;
    end

    reg [7:0] out309;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out309 = in0;
    end

    reg [7:0] out310;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out310 = in0;
    end

    reg [7:0] out311;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out311 = in0;
    end

    reg [7:0] out312;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out312 = in0;
    end

    reg [7:0] out313;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out313 = in0;
    end

    reg [7:0] out314;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out314 = in0;
    end

    reg [7:0] out315;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out315 = in0;
    end

    reg [7:0] out316;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out316 = in0;
    end

    reg [7:0] out317;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out317 = in0;
    end

    reg [7:0] out318;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out318 = in0;
    end

    reg [7:0] out319;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out319 = in0;
    end

    reg [7:0] out320;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out320 = in0;
    end

    reg [7:0] out321;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out321 = in0;
    end

    reg [7:0] out322;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out322 = in0;
    end

    reg [7:0] out323;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out323 = in0;
    end

    reg [7:0] out324;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out324 = in0;
    end

    reg [7:0] out325;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out325 = in0;
    end

    reg [7:0] out326;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out326 = in0;
    end

    reg [7:0] out327;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out327 = in0;
    end

    reg [7:0] out328;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out328 = in0;
    end

    reg [7:0] out329;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out329 = in0;
    end

    reg [7:0] out330;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out330 = in0;
    end

    reg [7:0] out331;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out331 = in0;
    end

    reg [7:0] out332;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out332 = in0;
    end

    reg [7:0] out333;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out333 = in0;
    end

    reg [7:0] out334;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out334 = in0;
    end

    reg [7:0] out335;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out335 = in0;
    end

    reg [7:0] out336;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out336 = in0;
    end

    reg [7:0] out337;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out337 = in0;
    end

    reg [7:0] out338;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out338 = in0;
    end

    reg [7:0] out339;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out339 = in0;
    end

    reg [7:0] out340;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out340 = in0;
    end

    reg [7:0] out341;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out341 = in0;
    end

    reg [7:0] out342;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out342 = in0;
    end

    reg [7:0] out343;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out343 = in0;
    end

    reg [7:0] out344;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out344 = in0;
    end

    reg [7:0] out345;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out345 = in0;
    end

    reg [7:0] out346;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out346 = in0;
    end

    reg [7:0] out347;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out347 = in0;
    end

    reg [7:0] out348;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out348 = in0;
    end

    reg [7:0] out349;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out349 = in0;
    end

    reg [7:0] out350;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out350 = in0;
    end

    reg [7:0] out351;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out351 = in0;
    end

    reg [7:0] out352;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out352 = in0;
    end

    reg [7:0] out353;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out353 = in0;
    end

    reg [7:0] out354;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out354 = in0;
    end

    reg [7:0] out355;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out355 = in0;
    end

    reg [7:0] out356;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out356 = in0;
    end

    reg [7:0] out357;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out357 = in0;
    end

    reg [7:0] out358;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out358 = in0;
    end

    reg [7:0] out359;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out359 = in0;
    end

    reg [7:0] out360;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out360 = in0;
    end

    reg [7:0] out361;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out361 = in0;
    end

    reg [7:0] out362;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out362 = in0;
    end

    reg [7:0] out363;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out363 = in0;
    end

    reg [7:0] out364;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out364 = in0;
    end

    reg [7:0] out365;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out365 = in0;
    end

    reg [7:0] out366;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out366 = in0;
    end

    reg [7:0] out367;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out367 = in0;
    end

    reg [7:0] out368;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out368 = in0;
    end

    reg [7:0] out369;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out369 = in0;
    end

    reg [7:0] out370;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out370 = in0;
    end

    reg [7:0] out371;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out371 = in0;
    end

    reg [7:0] out372;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out372 = in0;
    end

    reg [7:0] out373;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out373 = in0;
    end

    reg [7:0] out374;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out374 = in0;
    end

    reg [7:0] out375;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out375 = in0;
    end

    reg [7:0] out376;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out376 = in0;
    end

    reg [7:0] out377;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out377 = in0;
    end

    reg [7:0] out378;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out378 = in0;
    end

    reg [7:0] out379;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out379 = in0;
    end

    reg [7:0] out380;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out380 = in0;
    end

    reg [7:0] out381;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out381 = in0;
    end

    reg [7:0] out382;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out382 = in0;
    end

    reg [7:0] out383;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out383 = in0;
    end

    reg [7:0] out384;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out384 = in0;
    end

    reg [7:0] out385;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out385 = in0;
    end

    reg [7:0] out386;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out386 = in0;
    end

    reg [7:0] out387;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out387 = in0;
    end

    reg [7:0] out388;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out388 = in0;
    end

    reg [7:0] out389;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out389 = in0;
    end

    reg [7:0] out390;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out390 = in0;
    end

    reg [7:0] out391;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out391 = in0;
    end

    reg [7:0] out392;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out392 = in0;
    end

    reg [7:0] out393;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out393 = in0;
    end

    reg [7:0] out394;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out394 = in0;
    end

    reg [7:0] out395;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out395 = in0;
    end

    reg [7:0] out396;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out396 = in0;
    end

    reg [7:0] out397;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out397 = in0;
    end

    reg [7:0] out398;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out398 = in0;
    end

    reg [7:0] out399;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out399 = in0;
    end

    reg [7:0] out400;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out400 = in0;
    end

    reg [7:0] out401;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out401 = in0;
    end

    reg [7:0] out402;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out402 = in0;
    end

    reg [7:0] out403;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out403 = in0;
    end

    reg [7:0] out404;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out404 = in0;
    end

    reg [7:0] out405;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out405 = in0;
    end

    reg [7:0] out406;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out406 = in0;
    end

    reg [7:0] out407;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out407 = in0;
    end

    reg [7:0] out408;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out408 = in0;
    end

    reg [7:0] out409;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out409 = in0;
    end

    reg [7:0] out410;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out410 = in0;
    end

    reg [7:0] out411;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out411 = in0;
    end

    reg [7:0] out412;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out412 = in0;
    end

    reg [7:0] out413;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out413 = in0;
    end

    reg [7:0] out414;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out414 = in0;
    end

    reg [7:0] out415;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out415 = in0;
    end

    reg [7:0] out416;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out416 = in0;
    end

    reg [7:0] out417;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out417 = in0;
    end

    reg [7:0] out418;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out418 = in0;
    end

    reg [7:0] out419;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out419 = in0;
    end

    reg [7:0] out420;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out420 = in0;
    end

    reg [7:0] out421;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out421 = in0;
    end

    reg [7:0] out422;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out422 = in0;
    end

    reg [7:0] out423;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out423 = in0;
    end

    reg [7:0] out424;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out424 = in0;
    end

    reg [7:0] out425;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out425 = in0;
    end

    reg [7:0] out426;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out426 = in0;
    end

    reg [7:0] out427;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out427 = in0;
    end

    reg [7:0] out428;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out428 = in0;
    end

    reg [7:0] out429;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out429 = in0;
    end

    reg [7:0] out430;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out430 = in0;
    end

    reg [7:0] out431;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out431 = in0;
    end

    reg [7:0] out432;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out432 = in0;
    end

    reg [7:0] out433;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out433 = in0;
    end

    reg [7:0] out434;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out434 = in0;
    end

    reg [7:0] out435;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out435 = in0;
    end

    reg [7:0] out436;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out436 = in0;
    end

    reg [7:0] out437;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out437 = in0;
    end

    reg [7:0] out438;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out438 = in0;
    end

    reg [7:0] out439;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out439 = in0;
    end

    reg [7:0] out440;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out440 = in0;
    end

    reg [7:0] out441;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out441 = in0;
    end

    reg [7:0] out442;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out442 = in0;
    end

    reg [7:0] out443;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out443 = in0;
    end

    reg [7:0] out444;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out444 = in0;
    end

    reg [7:0] out445;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out445 = in0;
    end

    reg [7:0] out446;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out446 = in0;
    end

    reg [7:0] out447;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out447 = in0;
    end

    reg [7:0] out448;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out448 = in0;
    end

    reg [7:0] out449;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out449 = in0;
    end

    reg [7:0] out450;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out450 = in0;
    end

    reg [7:0] out451;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out451 = in0;
    end

    reg [7:0] out452;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out452 = in0;
    end

    reg [7:0] out453;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out453 = in0;
    end

    reg [7:0] out454;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out454 = in0;
    end

    reg [7:0] out455;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out455 = in0;
    end

    reg [7:0] out456;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out456 = in0;
    end

    reg [7:0] out457;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out457 = in0;
    end

    reg [7:0] out458;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out458 = in0;
    end

    reg [7:0] out459;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out459 = in0;
    end

    reg [7:0] out460;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out460 = in0;
    end

    reg [7:0] out461;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out461 = in0;
    end

    reg [7:0] out462;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out462 = in0;
    end

    reg [7:0] out463;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out463 = in0;
    end

    reg [7:0] out464;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out464 = in0;
    end

    reg [7:0] out465;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out465 = in0;
    end

    reg [7:0] out466;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out466 = in0;
    end

    reg [7:0] out467;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out467 = in0;
    end

    reg [7:0] out468;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out468 = in0;
    end

    reg [7:0] out469;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out469 = in0;
    end

    reg [7:0] out470;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out470 = in0;
    end

    reg [7:0] out471;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out471 = in0;
    end

    reg [7:0] out472;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out472 = in0;
    end

    reg [7:0] out473;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out473 = in0;
    end

    reg [7:0] out474;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out474 = in0;
    end

    reg [7:0] out475;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out475 = in0;
    end

    reg [7:0] out476;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out476 = in0;
    end

    reg [7:0] out477;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out477 = in0;
    end

    reg [7:0] out478;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out478 = in0;
    end

    reg [7:0] out479;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out479 = in0;
    end

    reg [7:0] out480;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out480 = in0;
    end

    reg [7:0] out481;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out481 = in0;
    end

    reg [7:0] out482;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out482 = in0;
    end

    reg [7:0] out483;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out483 = in0;
    end

    reg [7:0] out484;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out484 = in0;
    end

    reg [7:0] out485;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out485 = in0;
    end

    reg [7:0] out486;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out486 = in0;
    end

    reg [7:0] out487;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out487 = in0;
    end

    reg [7:0] out488;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out488 = in0;
    end

    reg [7:0] out489;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out489 = in0;
    end

    reg [7:0] out490;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out490 = in0;
    end

    reg [7:0] out491;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out491 = in0;
    end

    reg [7:0] out492;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out492 = in0;
    end

    reg [7:0] out493;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out493 = in0;
    end

    reg [7:0] out494;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out494 = in0;
    end

    reg [7:0] out495;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out495 = in0;
    end

    reg [7:0] out496;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out496 = in0;
    end

    reg [7:0] out497;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out497 = in0;
    end

    reg [7:0] out498;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out498 = in0;
    end

    reg [7:0] out499;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out499 = in0;
    end

    reg [7:0] out500;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out500 = in0;
    end

    reg [7:0] out501;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out501 = in0;
    end

    reg [7:0] out502;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out502 = in0;
    end

    reg [7:0] out503;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out503 = in0;
    end

    reg [7:0] out504;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out504 = in0;
    end

    reg [7:0] out505;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out505 = in0;
    end

    reg [7:0] out506;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out506 = in0;
    end

    reg [7:0] out507;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out507 = in0;
    end

    reg [7:0] out508;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out508 = in0;
    end

    reg [7:0] out509;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out509 = in0;
    end

    reg [7:0] out510;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out510 = in0;
    end

    reg [7:0] out511;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out511 = in0;
    end

    reg [7:0] out512;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out512 = in0;
    end

    reg [7:0] out513;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out513 = in0;
    end

    reg [7:0] out514;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out514 = in0;
    end

    reg [7:0] out515;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out515 = in0;
    end

    reg [7:0] out516;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out516 = in0;
    end

    reg [7:0] out517;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out517 = in0;
    end

    reg [7:0] out518;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out518 = in0;
    end

    reg [7:0] out519;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out519 = in0;
    end

    reg [7:0] out520;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out520 = in0;
    end

    reg [7:0] out521;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out521 = in0;
    end

    reg [7:0] out522;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out522 = in0;
    end

    reg [7:0] out523;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out523 = in0;
    end

    reg [7:0] out524;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out524 = in0;
    end

    reg [7:0] out525;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out525 = in0;
    end

    reg [7:0] out526;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out526 = in0;
    end

    reg [7:0] out527;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out527 = in0;
    end

    reg [7:0] out528;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out528 = in0;
    end

    reg [7:0] out529;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out529 = in0;
    end

    reg [7:0] out530;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out530 = in0;
    end

    reg [7:0] out531;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out531 = in0;
    end

    reg [7:0] out532;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out532 = in0;
    end

    reg [7:0] out533;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out533 = in0;
    end

    reg [7:0] out534;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out534 = in0;
    end

    reg [7:0] out535;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out535 = in0;
    end

    reg [7:0] out536;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out536 = in0;
    end

    reg [7:0] out537;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out537 = in0;
    end

    reg [7:0] out538;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out538 = in0;
    end

    reg [7:0] out539;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out539 = in0;
    end

    reg [7:0] out540;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out540 = in0;
    end

    reg [7:0] out541;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out541 = in0;
    end

    reg [7:0] out542;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out542 = in0;
    end

    reg [7:0] out543;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out543 = in0;
    end

    reg [7:0] out544;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out544 = in0;
    end

    reg [7:0] out545;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out545 = in0;
    end

    reg [7:0] out546;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out546 = in0;
    end

    reg [7:0] out547;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out547 = in0;
    end

    reg [7:0] out548;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out548 = in0;
    end

    reg [7:0] out549;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out549 = in0;
    end

    reg [7:0] out550;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out550 = in0;
    end

    reg [7:0] out551;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out551 = in0;
    end

    reg [7:0] out552;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out552 = in0;
    end

    reg [7:0] out553;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out553 = in0;
    end

    reg [7:0] out554;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out554 = in0;
    end

    reg [7:0] out555;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out555 = in0;
    end

    reg [7:0] out556;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out556 = in0;
    end

    reg [7:0] out557;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out557 = in0;
    end

    reg [7:0] out558;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out558 = in0;
    end

    reg [7:0] out559;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out559 = in0;
    end

    reg [7:0] out560;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out560 = in0;
    end

    reg [7:0] out561;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out561 = in0;
    end

    reg [7:0] out562;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out562 = in0;
    end

    reg [7:0] out563;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out563 = in0;
    end

    reg [7:0] out564;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out564 = in0;
    end

    reg [7:0] out565;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out565 = in0;
    end

    reg [7:0] out566;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out566 = in0;
    end

    reg [7:0] out567;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out567 = in0;
    end

    reg [7:0] out568;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out568 = in0;
    end

    reg [7:0] out569;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out569 = in0;
    end

    reg [7:0] out570;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out570 = in0;
    end

    reg [7:0] out571;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out571 = in0;
    end

    reg [7:0] out572;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out572 = in0;
    end

    reg [7:0] out573;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out573 = in0;
    end

    reg [7:0] out574;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out574 = in0;
    end

    reg [7:0] out575;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out575 = in0;
    end

    reg [7:0] out576;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out576 = in0;
    end

    reg [7:0] out577;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out577 = in0;
    end

    reg [7:0] out578;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out578 = in0;
    end

    reg [7:0] out579;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out579 = in0;
    end

    reg [7:0] out580;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out580 = in0;
    end

    reg [7:0] out581;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out581 = in0;
    end

    reg [7:0] out582;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out582 = in0;
    end

    reg [7:0] out583;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out583 = in0;
    end

    reg [7:0] out584;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out584 = in0;
    end

    reg [7:0] out585;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out585 = in0;
    end

    reg [7:0] out586;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out586 = in0;
    end

    reg [7:0] out587;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out587 = in0;
    end

    reg [7:0] out588;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out588 = in0;
    end

    reg [7:0] out589;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out589 = in0;
    end

    reg [7:0] out590;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out590 = in0;
    end

    reg [7:0] out591;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out591 = in0;
    end

    reg [7:0] out592;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out592 = in0;
    end

    reg [7:0] out593;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out593 = in0;
    end

    reg [7:0] out594;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out594 = in0;
    end

    reg [7:0] out595;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out595 = in0;
    end

    reg [7:0] out596;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out596 = in0;
    end

    reg [7:0] out597;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out597 = in0;
    end

    reg [7:0] out598;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out598 = in0;
    end

    reg [7:0] out599;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out599 = in0;
    end

    reg [7:0] out600;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out600 = in0;
    end

    reg [7:0] out601;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out601 = in0;
    end

    reg [7:0] out602;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out602 = in0;
    end

    reg [7:0] out603;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out603 = in0;
    end

    reg [7:0] out604;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out604 = in0;
    end

    reg [7:0] out605;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out605 = in0;
    end

    reg [7:0] out606;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out606 = in0;
    end

    reg [7:0] out607;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out607 = in0;
    end

    reg [7:0] out608;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out608 = in0;
    end

    reg [7:0] out609;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out609 = in0;
    end

    reg [7:0] out610;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out610 = in0;
    end

    reg [7:0] out611;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out611 = in0;
    end

    reg [7:0] out612;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out612 = in0;
    end

    reg [7:0] out613;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out613 = in0;
    end

    reg [7:0] out614;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out614 = in0;
    end

    reg [7:0] out615;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out615 = in0;
    end

    reg [7:0] out616;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out616 = in0;
    end

    reg [7:0] out617;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out617 = in0;
    end

    reg [7:0] out618;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out618 = in0;
    end

    reg [7:0] out619;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out619 = in0;
    end

    reg [7:0] out620;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out620 = in0;
    end

    reg [7:0] out621;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out621 = in0;
    end

    reg [7:0] out622;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out622 = in0;
    end

    reg [7:0] out623;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out623 = in0;
    end

    reg [7:0] out624;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out624 = in0;
    end

    reg [7:0] out625;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out625 = in0;
    end

    reg [7:0] out626;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out626 = in0;
    end

    reg [7:0] out627;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out627 = in0;
    end

    reg [7:0] out628;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out628 = in0;
    end

    reg [7:0] out629;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out629 = in0;
    end

    reg [7:0] out630;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out630 = in0;
    end

    reg [7:0] out631;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out631 = in0;
    end

    reg [7:0] out632;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out632 = in0;
    end

    reg [7:0] out633;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out633 = in0;
    end

    reg [7:0] out634;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out634 = in0;
    end

    reg [7:0] out635;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out635 = in0;
    end

    reg [7:0] out636;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out636 = in0;
    end

    reg [7:0] out637;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out637 = in0;
    end

    reg [7:0] out638;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out638 = in0;
    end

    reg [7:0] out639;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out639 = in0;
    end

    reg [7:0] out640;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out640 = in0;
    end

    reg [7:0] out641;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out641 = in0;
    end

    reg [7:0] out642;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out642 = in0;
    end

    reg [7:0] out643;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out643 = in0;
    end

    reg [7:0] out644;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out644 = in0;
    end

    reg [7:0] out645;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out645 = in0;
    end

    reg [7:0] out646;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out646 = in0;
    end

    reg [7:0] out647;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out647 = in0;
    end

    reg [7:0] out648;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out648 = in0;
    end

    reg [7:0] out649;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out649 = in0;
    end

    reg [7:0] out650;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out650 = in0;
    end

    reg [7:0] out651;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out651 = in0;
    end

    reg [7:0] out652;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out652 = in0;
    end

    reg [7:0] out653;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out653 = in0;
    end

    reg [7:0] out654;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out654 = in0;
    end

    reg [7:0] out655;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out655 = in0;
    end

    reg [7:0] out656;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out656 = in0;
    end

    reg [7:0] out657;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out657 = in0;
    end

    reg [7:0] out658;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out658 = in0;
    end

    reg [7:0] out659;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out659 = in0;
    end

    reg [7:0] out660;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out660 = in0;
    end

    reg [7:0] out661;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out661 = in0;
    end

    reg [7:0] out662;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out662 = in0;
    end

    reg [7:0] out663;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out663 = in0;
    end

    reg [7:0] out664;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out664 = in0;
    end

    reg [7:0] out665;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out665 = in0;
    end

    reg [7:0] out666;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out666 = in0;
    end

    reg [7:0] out667;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out667 = in0;
    end

    reg [7:0] out668;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out668 = in0;
    end

    reg [7:0] out669;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out669 = in0;
    end

    reg [7:0] out670;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out670 = in0;
    end

    reg [7:0] out671;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out671 = in0;
    end

    reg [7:0] out672;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out672 = in0;
    end

    reg [7:0] out673;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out673 = in0;
    end

    reg [7:0] out674;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out674 = in0;
    end

    reg [7:0] out675;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out675 = in0;
    end

    reg [7:0] out676;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out676 = in0;
    end

    reg [7:0] out677;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out677 = in0;
    end

    reg [7:0] out678;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out678 = in0;
    end

    reg [7:0] out679;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out679 = in0;
    end

    reg [7:0] out680;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out680 = in0;
    end

    reg [7:0] out681;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out681 = in0;
    end

    reg [7:0] out682;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out682 = in0;
    end

    reg [7:0] out683;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out683 = in0;
    end

    reg [7:0] out684;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out684 = in0;
    end

    reg [7:0] out685;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out685 = in0;
    end

    reg [7:0] out686;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out686 = in0;
    end

    reg [7:0] out687;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out687 = in0;
    end

    reg [7:0] out688;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out688 = in0;
    end

    reg [7:0] out689;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out689 = in0;
    end

    reg [7:0] out690;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out690 = in0;
    end

    reg [7:0] out691;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out691 = in0;
    end

    reg [7:0] out692;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out692 = in0;
    end

    reg [7:0] out693;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out693 = in0;
    end

    reg [7:0] out694;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out694 = in0;
    end

    reg [7:0] out695;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out695 = in0;
    end

    reg [7:0] out696;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out696 = in0;
    end

    reg [7:0] out697;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out697 = in0;
    end

    reg [7:0] out698;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out698 = in0;
    end

    reg [7:0] out699;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out699 = in0;
    end

    reg [7:0] out700;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out700 = in0;
    end

    reg [7:0] out701;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out701 = in0;
    end

    reg [7:0] out702;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out702 = in0;
    end

    reg [7:0] out703;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out703 = in0;
    end

    reg [7:0] out704;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out704 = in0;
    end

    reg [7:0] out705;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out705 = in0;
    end

    reg [7:0] out706;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out706 = in0;
    end

    reg [7:0] out707;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out707 = in0;
    end

    reg [7:0] out708;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out708 = in0;
    end

    reg [7:0] out709;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out709 = in0;
    end

    reg [7:0] out710;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out710 = in0;
    end

    reg [7:0] out711;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out711 = in0;
    end

    reg [7:0] out712;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out712 = in0;
    end

    reg [7:0] out713;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out713 = in0;
    end

    reg [7:0] out714;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out714 = in0;
    end

    reg [7:0] out715;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out715 = in0;
    end

    reg [7:0] out716;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out716 = in0;
    end

    reg [7:0] out717;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out717 = in0;
    end

    reg [7:0] out718;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out718 = in0;
    end

    reg [7:0] out719;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out719 = in0;
    end

    reg [7:0] out720;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out720 = in0;
    end

    reg [7:0] out721;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out721 = in0;
    end

    reg [7:0] out722;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out722 = in0;
    end

    reg [7:0] out723;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out723 = in0;
    end

    reg [7:0] out724;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out724 = in0;
    end

    reg [7:0] out725;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out725 = in0;
    end

    reg [7:0] out726;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out726 = in0;
    end

    reg [7:0] out727;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out727 = in0;
    end

    reg [7:0] out728;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out728 = in0;
    end

    reg [7:0] out729;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out729 = in0;
    end

    reg [7:0] out730;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out730 = in0;
    end

    reg [7:0] out731;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out731 = in0;
    end

    reg [7:0] out732;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out732 = in0;
    end

    reg [7:0] out733;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out733 = in0;
    end

    reg [7:0] out734;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out734 = in0;
    end

    reg [7:0] out735;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out735 = in0;
    end

    reg [7:0] out736;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out736 = in0;
    end

    reg [7:0] out737;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out737 = in0;
    end

    reg [7:0] out738;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out738 = in0;
    end

    reg [7:0] out739;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out739 = in0;
    end

    reg [7:0] out740;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out740 = in0;
    end

    reg [7:0] out741;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out741 = in0;
    end

    reg [7:0] out742;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out742 = in0;
    end

    reg [7:0] out743;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out743 = in0;
    end

    reg [7:0] out744;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out744 = in0;
    end

    reg [7:0] out745;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out745 = in0;
    end

    reg [7:0] out746;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out746 = in0;
    end

    reg [7:0] out747;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out747 = in0;
    end

    reg [7:0] out748;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out748 = in0;
    end

    reg [7:0] out749;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out749 = in0;
    end

    reg [7:0] out750;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out750 = in0;
    end

    reg [7:0] out751;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out751 = in0;
    end

    reg [7:0] out752;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out752 = in0;
    end

    reg [7:0] out753;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out753 = in0;
    end

    reg [7:0] out754;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out754 = in0;
    end

    reg [7:0] out755;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out755 = in0;
    end

    reg [7:0] out756;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out756 = in0;
    end

    reg [7:0] out757;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out757 = in0;
    end

    reg [7:0] out758;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out758 = in0;
    end

    reg [7:0] out759;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out759 = in0;
    end

    reg [7:0] out760;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out760 = in0;
    end

    reg [7:0] out761;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out761 = in0;
    end

    reg [7:0] out762;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out762 = in0;
    end

    reg [7:0] out763;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out763 = in0;
    end

    reg [7:0] out764;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out764 = in0;
    end

    reg [7:0] out765;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out765 = in0;
    end

    reg [7:0] out766;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out766 = in0;
    end

    reg [7:0] out767;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out767 = in0;
    end

    reg [7:0] out768;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out768 = in0;
    end

    reg [7:0] out769;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out769 = in0;
    end

    reg [7:0] out770;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out770 = in0;
    end

    reg [7:0] out771;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out771 = in0;
    end

    reg [7:0] out772;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out772 = in0;
    end

    reg [7:0] out773;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out773 = in0;
    end

    reg [7:0] out774;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out774 = in0;
    end

    reg [7:0] out775;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out775 = in0;
    end

    reg [7:0] out776;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out776 = in0;
    end

    reg [7:0] out777;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out777 = in0;
    end

    reg [7:0] out778;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out778 = in0;
    end

    reg [7:0] out779;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out779 = in0;
    end

    reg [7:0] out780;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out780 = in0;
    end

    reg [7:0] out781;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out781 = in0;
    end

    reg [7:0] out782;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out782 = in0;
    end

    reg [7:0] out783;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out783 = in0;
    end

    reg [7:0] out784;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out784 = in0;
    end

    reg [7:0] out785;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out785 = in0;
    end

    reg [7:0] out786;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out786 = in0;
    end

    reg [7:0] out787;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out787 = in0;
    end

    reg [7:0] out788;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out788 = in0;
    end

    reg [7:0] out789;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out789 = in0;
    end

    reg [7:0] out790;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out790 = in0;
    end

    reg [7:0] out791;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out791 = in0;
    end

    reg [7:0] out792;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out792 = in0;
    end

    reg [7:0] out793;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out793 = in0;
    end

    reg [7:0] out794;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out794 = in0;
    end

    reg [7:0] out795;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out795 = in0;
    end

    reg [7:0] out796;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out796 = in0;
    end

    reg [7:0] out797;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out797 = in0;
    end

    reg [7:0] out798;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out798 = in0;
    end

    reg [7:0] out799;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out799 = in0;
    end

    reg [7:0] out800;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out800 = in0;
    end

    reg [7:0] out801;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out801 = in0;
    end

    reg [7:0] out802;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out802 = in0;
    end

    reg [7:0] out803;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out803 = in0;
    end

    reg [7:0] out804;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out804 = in0;
    end

    reg [7:0] out805;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out805 = in0;
    end

    reg [7:0] out806;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out806 = in0;
    end

    reg [7:0] out807;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out807 = in0;
    end

    reg [7:0] out808;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out808 = in0;
    end

    reg [7:0] out809;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out809 = in0;
    end

    reg [7:0] out810;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out810 = in0;
    end

    reg [7:0] out811;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out811 = in0;
    end

    reg [7:0] out812;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out812 = in0;
    end

    reg [7:0] out813;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out813 = in0;
    end

    reg [7:0] out814;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out814 = in0;
    end

    reg [7:0] out815;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out815 = in0;
    end

    reg [7:0] out816;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out816 = in0;
    end

    reg [7:0] out817;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out817 = in0;
    end

    reg [7:0] out818;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out818 = in0;
    end

    reg [7:0] out819;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out819 = in0;
    end

    reg [7:0] out820;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out820 = in0;
    end

    reg [7:0] out821;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out821 = in0;
    end

    reg [7:0] out822;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out822 = in0;
    end

    reg [7:0] out823;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out823 = in0;
    end

    reg [7:0] out824;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out824 = in0;
    end

    reg [7:0] out825;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out825 = in0;
    end

    reg [7:0] out826;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out826 = in0;
    end

    reg [7:0] out827;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out827 = in0;
    end

    reg [7:0] out828;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out828 = in0;
    end

    reg [7:0] out829;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out829 = in0;
    end

    reg [7:0] out830;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out830 = in0;
    end

    reg [7:0] out831;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out831 = in0;
    end

    reg [7:0] out832;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out832 = in0;
    end

    reg [7:0] out833;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out833 = in0;
    end

    reg [7:0] out834;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out834 = in0;
    end

    reg [7:0] out835;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out835 = in0;
    end

    reg [7:0] out836;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out836 = in0;
    end

    reg [7:0] out837;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out837 = in0;
    end

    reg [7:0] out838;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out838 = in0;
    end

    reg [7:0] out839;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out839 = in0;
    end

    reg [7:0] out840;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out840 = in0;
    end

    reg [7:0] out841;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out841 = in0;
    end

    reg [7:0] out842;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out842 = in0;
    end

    reg [7:0] out843;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out843 = in0;
    end

    reg [7:0] out844;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out844 = in0;
    end

    reg [7:0] out845;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out845 = in0;
    end

    reg [7:0] out846;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out846 = in0;
    end

    reg [7:0] out847;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out847 = in0;
    end

    reg [7:0] out848;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out848 = in0;
    end

    reg [7:0] out849;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out849 = in0;
    end

    reg [7:0] out850;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out850 = in0;
    end

    reg [7:0] out851;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out851 = in0;
    end

    reg [7:0] out852;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out852 = in0;
    end

    reg [7:0] out853;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out853 = in0;
    end

    reg [7:0] out854;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out854 = in0;
    end

    reg [7:0] out855;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out855 = in0;
    end

    reg [7:0] out856;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out856 = in0;
    end

    reg [7:0] out857;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out857 = in0;
    end

    reg [7:0] out858;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out858 = in0;
    end

    reg [7:0] out859;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out859 = in0;
    end

    reg [7:0] out860;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out860 = in0;
    end

    reg [7:0] out861;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out861 = in0;
    end

    reg [7:0] out862;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out862 = in0;
    end

    reg [7:0] out863;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out863 = in0;
    end

    reg [7:0] out864;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out864 = in0;
    end

    reg [7:0] out865;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out865 = in0;
    end

    reg [7:0] out866;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out866 = in0;
    end

    reg [7:0] out867;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out867 = in0;
    end

    reg [7:0] out868;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out868 = in0;
    end

    reg [7:0] out869;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out869 = in0;
    end

    reg [7:0] out870;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out870 = in0;
    end

    reg [7:0] out871;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out871 = in0;
    end

    reg [7:0] out872;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out872 = in0;
    end

    reg [7:0] out873;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out873 = in0;
    end

    reg [7:0] out874;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out874 = in0;
    end

    reg [7:0] out875;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out875 = in0;
    end

    reg [7:0] out876;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out876 = in0;
    end

    reg [7:0] out877;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out877 = in0;
    end

    reg [7:0] out878;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out878 = in0;
    end

    reg [7:0] out879;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out879 = in0;
    end

    reg [7:0] out880;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out880 = in0;
    end

    reg [7:0] out881;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out881 = in0;
    end

    reg [7:0] out882;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out882 = in0;
    end

    reg [7:0] out883;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out883 = in0;
    end

    reg [7:0] out884;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out884 = in0;
    end

    reg [7:0] out885;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out885 = in0;
    end

    reg [7:0] out886;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out886 = in0;
    end

    reg [7:0] out887;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out887 = in0;
    end

    reg [7:0] out888;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out888 = in0;
    end

    reg [7:0] out889;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out889 = in0;
    end

    reg [7:0] out890;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out890 = in0;
    end

    reg [7:0] out891;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out891 = in0;
    end

    reg [7:0] out892;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out892 = in0;
    end

    reg [7:0] out893;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out893 = in0;
    end

    reg [7:0] out894;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out894 = in0;
    end

    reg [7:0] out895;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out895 = in0;
    end

    reg [7:0] out896;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out896 = in0;
    end

    reg [7:0] out897;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out897 = in0;
    end

    reg [7:0] out898;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out898 = in0;
    end

    reg [7:0] out899;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out899 = in0;
    end

    reg [7:0] out900;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out900 = in0;
    end

    reg [7:0] out901;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out901 = in0;
    end

    reg [7:0] out902;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out902 = in0;
    end

    reg [7:0] out903;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out903 = in0;
    end

    reg [7:0] out904;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out904 = in0;
    end

    reg [7:0] out905;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out905 = in0;
    end

    reg [7:0] out906;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out906 = in0;
    end

    reg [7:0] out907;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out907 = in0;
    end

    reg [7:0] out908;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out908 = in0;
    end

    reg [7:0] out909;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out909 = in0;
    end

    reg [7:0] out910;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out910 = in0;
    end

    reg [7:0] out911;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out911 = in0;
    end

    reg [7:0] out912;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out912 = in0;
    end

    reg [7:0] out913;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out913 = in0;
    end

    reg [7:0] out914;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out914 = in0;
    end

    reg [7:0] out915;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out915 = in0;
    end

    reg [7:0] out916;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out916 = in0;
    end

    reg [7:0] out917;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out917 = in0;
    end

    reg [7:0] out918;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out918 = in0;
    end

    reg [7:0] out919;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out919 = in0;
    end

    reg [7:0] out920;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out920 = in0;
    end

    reg [7:0] out921;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out921 = in0;
    end

    reg [7:0] out922;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out922 = in0;
    end

    reg [7:0] out923;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out923 = in0;
    end

    reg [7:0] out924;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out924 = in0;
    end

    reg [7:0] out925;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out925 = in0;
    end

    reg [7:0] out926;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out926 = in0;
    end

    reg [7:0] out927;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out927 = in0;
    end

    reg [7:0] out928;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out928 = in0;
    end

    reg [7:0] out929;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out929 = in0;
    end

    reg [7:0] out930;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out930 = in0;
    end

    reg [7:0] out931;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out931 = in0;
    end

    reg [7:0] out932;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out932 = in0;
    end

    reg [7:0] out933;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out933 = in0;
    end

    reg [7:0] out934;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out934 = in0;
    end

    reg [7:0] out935;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out935 = in0;
    end

    reg [7:0] out936;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out936 = in0;
    end

    reg [7:0] out937;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out937 = in0;
    end

    reg [7:0] out938;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out938 = in0;
    end

    reg [7:0] out939;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out939 = in0;
    end

    reg [7:0] out940;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out940 = in0;
    end

    reg [7:0] out941;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out941 = in0;
    end

    reg [7:0] out942;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out942 = in0;
    end

    reg [7:0] out943;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out943 = in0;
    end

    reg [7:0] out944;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out944 = in0;
    end

    reg [7:0] out945;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out945 = in0;
    end

    reg [7:0] out946;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out946 = in0;
    end

    reg [7:0] out947;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out947 = in0;
    end

    reg [7:0] out948;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out948 = in0;
    end

    reg [7:0] out949;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out949 = in0;
    end

    reg [7:0] out950;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out950 = in0;
    end

    reg [7:0] out951;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out951 = in0;
    end

    reg [7:0] out952;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out952 = in0;
    end

    reg [7:0] out953;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out953 = in0;
    end

    reg [7:0] out954;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out954 = in0;
    end

    reg [7:0] out955;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out955 = in0;
    end

    reg [7:0] out956;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out956 = in0;
    end

    reg [7:0] out957;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out957 = in0;
    end

    reg [7:0] out958;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out958 = in0;
    end

    reg [7:0] out959;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out959 = in0;
    end

    reg [7:0] out960;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out960 = in0;
    end

    reg [7:0] out961;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out961 = in0;
    end

    reg [7:0] out962;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out962 = in0;
    end

    reg [7:0] out963;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out963 = in0;
    end

    reg [7:0] out964;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out964 = in0;
    end

    reg [7:0] out965;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out965 = in0;
    end

    reg [7:0] out966;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out966 = in0;
    end

    reg [7:0] out967;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out967 = in0;
    end

    reg [7:0] out968;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out968 = in0;
    end

    reg [7:0] out969;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out969 = in0;
    end

    reg [7:0] out970;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out970 = in0;
    end

    reg [7:0] out971;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out971 = in0;
    end

    reg [7:0] out972;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out972 = in0;
    end

    reg [7:0] out973;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out973 = in0;
    end

    reg [7:0] out974;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out974 = in0;
    end

    reg [7:0] out975;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out975 = in0;
    end

    reg [7:0] out976;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out976 = in0;
    end

    reg [7:0] out977;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out977 = in0;
    end

    reg [7:0] out978;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out978 = in0;
    end

    reg [7:0] out979;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out979 = in0;
    end

    reg [7:0] out980;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out980 = in0;
    end

    reg [7:0] out981;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out981 = in0;
    end

    reg [7:0] out982;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out982 = in0;
    end

    reg [7:0] out983;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out983 = in0;
    end

    reg [7:0] out984;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out984 = in0;
    end

    reg [7:0] out985;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out985 = in0;
    end

    reg [7:0] out986;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out986 = in0;
    end

    reg [7:0] out987;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out987 = in0;
    end

    reg [7:0] out988;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out988 = in0;
    end

    reg [7:0] out989;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out989 = in0;
    end

    reg [7:0] out990;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out990 = in0;
    end

    reg [7:0] out991;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out991 = in0;
    end

    reg [7:0] out992;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out992 = in0;
    end

    reg [7:0] out993;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out993 = in0;
    end

    reg [7:0] out994;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out994 = in0;
    end

    reg [7:0] out995;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out995 = in0;
    end

    reg [7:0] out996;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out996 = in0;
    end

    reg [7:0] out997;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out997 = in0;
    end

    reg [7:0] out998;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out998 = in0;
    end

    reg [7:0] out999;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out999 = in0;
    end

    reg [7:0] out1000;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1000 = in0;
    end

    reg [7:0] out1001;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1001 = in0;
    end

    reg [7:0] out1002;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1002 = in0;
    end

    reg [7:0] out1003;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1003 = in0;
    end

    reg [7:0] out1004;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1004 = in0;
    end

    reg [7:0] out1005;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1005 = in0;
    end

    reg [7:0] out1006;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1006 = in0;
    end

    reg [7:0] out1007;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1007 = in0;
    end

    reg [7:0] out1008;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1008 = in0;
    end

    reg [7:0] out1009;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1009 = in0;
    end

    reg [7:0] out1010;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1010 = in0;
    end

    reg [7:0] out1011;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1011 = in0;
    end

    reg [7:0] out1012;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1012 = in0;
    end

    reg [7:0] out1013;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1013 = in0;
    end

    reg [7:0] out1014;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1014 = in0;
    end

    reg [7:0] out1015;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1015 = in0;
    end

    reg [7:0] out1016;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1016 = in0;
    end

    reg [7:0] out1017;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1017 = in0;
    end

    reg [7:0] out1018;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1018 = in0;
    end

    reg [7:0] out1019;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1019 = in0;
    end

    reg [7:0] out1020;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1020 = in0;
    end

    reg [7:0] out1021;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1021 = in0;
    end

    reg [7:0] out1022;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1022 = in0;
    end

    reg [7:0] out1023;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1023 = in0;
    end

    reg [7:0] out1024;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1024 = in0;
    end

    reg [7:0] out1025;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1025 = in0;
    end

    reg [7:0] out1026;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1026 = in0;
    end

    reg [7:0] out1027;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1027 = in0;
    end

    reg [7:0] out1028;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1028 = in0;
    end

    reg [7:0] out1029;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1029 = in0;
    end

    reg [7:0] out1030;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1030 = in0;
    end

    reg [7:0] out1031;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1031 = in0;
    end

    reg [7:0] out1032;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1032 = in0;
    end

    reg [7:0] out1033;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1033 = in0;
    end

    reg [7:0] out1034;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1034 = in0;
    end

    reg [7:0] out1035;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1035 = in0;
    end

    reg [7:0] out1036;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1036 = in0;
    end

    reg [7:0] out1037;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1037 = in0;
    end

    reg [7:0] out1038;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1038 = in0;
    end

    reg [7:0] out1039;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1039 = in0;
    end

    reg [7:0] out1040;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1040 = in0;
    end

    reg [7:0] out1041;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1041 = in0;
    end

    reg [7:0] out1042;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1042 = in0;
    end

    reg [7:0] out1043;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1043 = in0;
    end

    reg [7:0] out1044;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1044 = in0;
    end

    reg [7:0] out1045;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1045 = in0;
    end

    reg [7:0] out1046;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1046 = in0;
    end

    reg [7:0] out1047;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1047 = in0;
    end

    reg [7:0] out1048;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1048 = in0;
    end

    reg [7:0] out1049;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1049 = in0;
    end

    reg [7:0] out1050;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1050 = in0;
    end

    reg [7:0] out1051;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1051 = in0;
    end

    reg [7:0] out1052;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1052 = in0;
    end

    reg [7:0] out1053;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1053 = in0;
    end

    reg [7:0] out1054;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1054 = in0;
    end

    reg [7:0] out1055;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1055 = in0;
    end

    reg [7:0] out1056;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1056 = in0;
    end

    reg [7:0] out1057;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1057 = in0;
    end

    reg [7:0] out1058;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1058 = in0;
    end

    reg [7:0] out1059;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1059 = in0;
    end

    reg [7:0] out1060;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1060 = in0;
    end

    reg [7:0] out1061;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1061 = in0;
    end

    reg [7:0] out1062;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1062 = in0;
    end

    reg [7:0] out1063;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1063 = in0;
    end

    reg [7:0] out1064;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1064 = in0;
    end

    reg [7:0] out1065;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1065 = in0;
    end

    reg [7:0] out1066;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1066 = in0;
    end

    reg [7:0] out1067;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1067 = in0;
    end

    reg [7:0] out1068;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1068 = in0;
    end

    reg [7:0] out1069;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1069 = in0;
    end

    reg [7:0] out1070;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1070 = in0;
    end

    reg [7:0] out1071;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1071 = in0;
    end

    reg [7:0] out1072;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1072 = in0;
    end

    reg [7:0] out1073;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1073 = in0;
    end

    reg [7:0] out1074;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1074 = in0;
    end

    reg [7:0] out1075;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1075 = in0;
    end

    reg [7:0] out1076;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1076 = in0;
    end

    reg [7:0] out1077;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1077 = in0;
    end

    reg [7:0] out1078;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1078 = in0;
    end

    reg [7:0] out1079;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1079 = in0;
    end

    reg [7:0] out1080;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1080 = in0;
    end

    reg [7:0] out1081;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1081 = in0;
    end

    reg [7:0] out1082;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1082 = in0;
    end

    reg [7:0] out1083;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1083 = in0;
    end

    reg [7:0] out1084;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1084 = in0;
    end

    reg [7:0] out1085;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1085 = in0;
    end

    reg [7:0] out1086;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1086 = in0;
    end

    reg [7:0] out1087;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1087 = in0;
    end

    reg [7:0] out1088;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1088 = in0;
    end

    reg [7:0] out1089;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1089 = in0;
    end

    reg [7:0] out1090;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1090 = in0;
    end

    reg [7:0] out1091;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1091 = in0;
    end

    reg [7:0] out1092;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1092 = in0;
    end

    reg [7:0] out1093;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1093 = in0;
    end

    reg [7:0] out1094;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1094 = in0;
    end

    reg [7:0] out1095;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1095 = in0;
    end

    reg [7:0] out1096;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1096 = in0;
    end

    reg [7:0] out1097;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1097 = in0;
    end

    reg [7:0] out1098;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1098 = in0;
    end

    reg [7:0] out1099;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1099 = in0;
    end

    reg [7:0] out1100;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1100 = in0;
    end

    reg [7:0] out1101;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1101 = in0;
    end

    reg [7:0] out1102;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1102 = in0;
    end

    reg [7:0] out1103;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1103 = in0;
    end

    reg [7:0] out1104;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1104 = in0;
    end

    reg [7:0] out1105;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1105 = in0;
    end

    reg [7:0] out1106;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1106 = in0;
    end

    reg [7:0] out1107;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1107 = in0;
    end

    reg [7:0] out1108;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1108 = in0;
    end

    reg [7:0] out1109;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1109 = in0;
    end

    reg [7:0] out1110;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1110 = in0;
    end

    reg [7:0] out1111;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1111 = in0;
    end

    reg [7:0] out1112;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1112 = in0;
    end

    reg [7:0] out1113;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1113 = in0;
    end

    reg [7:0] out1114;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1114 = in0;
    end

    reg [7:0] out1115;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1115 = in0;
    end

    reg [7:0] out1116;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1116 = in0;
    end

    reg [7:0] out1117;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1117 = in0;
    end

    reg [7:0] out1118;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1118 = in0;
    end

    reg [7:0] out1119;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1119 = in0;
    end

    reg [7:0] out1120;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1120 = in0;
    end

    reg [7:0] out1121;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1121 = in0;
    end

    reg [7:0] out1122;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1122 = in0;
    end

    reg [7:0] out1123;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1123 = in0;
    end

    reg [7:0] out1124;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1124 = in0;
    end

    reg [7:0] out1125;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1125 = in0;
    end

    reg [7:0] out1126;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1126 = in0;
    end

    reg [7:0] out1127;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1127 = in0;
    end

    reg [7:0] out1128;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1128 = in0;
    end

    reg [7:0] out1129;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1129 = in0;
    end

    reg [7:0] out1130;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1130 = in0;
    end

    reg [7:0] out1131;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1131 = in0;
    end

    reg [7:0] out1132;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1132 = in0;
    end

    reg [7:0] out1133;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1133 = in0;
    end

    reg [7:0] out1134;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1134 = in0;
    end

    reg [7:0] out1135;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1135 = in0;
    end

    reg [7:0] out1136;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1136 = in0;
    end

    reg [7:0] out1137;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1137 = in0;
    end

    reg [7:0] out1138;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1138 = in0;
    end

    reg [7:0] out1139;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1139 = in0;
    end

    reg [7:0] out1140;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1140 = in0;
    end

    reg [7:0] out1141;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1141 = in0;
    end

    reg [7:0] out1142;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1142 = in0;
    end

    reg [7:0] out1143;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1143 = in0;
    end

    reg [7:0] out1144;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1144 = in0;
    end

    reg [7:0] out1145;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1145 = in0;
    end

    reg [7:0] out1146;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1146 = in0;
    end

    reg [7:0] out1147;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1147 = in0;
    end

    reg [7:0] out1148;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1148 = in0;
    end

    reg [7:0] out1149;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1149 = in0;
    end

    reg [7:0] out1150;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1150 = in0;
    end

    reg [7:0] out1151;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1151 = in0;
    end

    reg [7:0] out1152;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1152 = in0;
    end

    reg [7:0] out1153;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1153 = in0;
    end

    reg [7:0] out1154;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1154 = in0;
    end

    reg [7:0] out1155;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1155 = in0;
    end

    reg [7:0] out1156;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1156 = in0;
    end

    reg [7:0] out1157;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1157 = in0;
    end

    reg [7:0] out1158;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1158 = in0;
    end

    reg [7:0] out1159;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1159 = in0;
    end

    reg [7:0] out1160;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1160 = in0;
    end

    reg [7:0] out1161;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1161 = in0;
    end

    reg [7:0] out1162;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1162 = in0;
    end

    reg [7:0] out1163;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1163 = in0;
    end

    reg [7:0] out1164;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1164 = in0;
    end

    reg [7:0] out1165;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1165 = in0;
    end

    reg [7:0] out1166;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1166 = in0;
    end

    reg [7:0] out1167;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1167 = in0;
    end

    reg [7:0] out1168;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1168 = in0;
    end

    reg [7:0] out1169;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1169 = in0;
    end

    reg [7:0] out1170;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1170 = in0;
    end

    reg [7:0] out1171;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1171 = in0;
    end

    reg [7:0] out1172;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1172 = in0;
    end

    reg [7:0] out1173;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1173 = in0;
    end

    reg [7:0] out1174;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1174 = in0;
    end

    reg [7:0] out1175;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1175 = in0;
    end

    reg [7:0] out1176;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1176 = in0;
    end

    reg [7:0] out1177;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1177 = in0;
    end

    reg [7:0] out1178;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1178 = in0;
    end

    reg [7:0] out1179;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1179 = in0;
    end

    reg [7:0] out1180;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1180 = in0;
    end

    reg [7:0] out1181;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1181 = in0;
    end

    reg [7:0] out1182;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1182 = in0;
    end

    reg [7:0] out1183;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1183 = in0;
    end

    reg [7:0] out1184;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1184 = in0;
    end

    reg [7:0] out1185;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1185 = in0;
    end

    reg [7:0] out1186;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1186 = in0;
    end

    reg [7:0] out1187;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1187 = in0;
    end

    reg [7:0] out1188;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1188 = in0;
    end

    reg [7:0] out1189;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1189 = in0;
    end

    reg [7:0] out1190;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1190 = in0;
    end

    reg [7:0] out1191;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1191 = in0;
    end

    reg [7:0] out1192;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1192 = in0;
    end

    reg [7:0] out1193;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1193 = in0;
    end

    reg [7:0] out1194;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1194 = in0;
    end

    reg [7:0] out1195;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1195 = in0;
    end

    reg [7:0] out1196;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1196 = in0;
    end

    reg [7:0] out1197;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1197 = in0;
    end

    reg [7:0] out1198;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1198 = in0;
    end

    reg [7:0] out1199;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1199 = in0;
    end

    reg [7:0] out1200;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1200 = in0;
    end

    reg [7:0] out1201;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1201 = in0;
    end

    reg [7:0] out1202;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1202 = in0;
    end

    reg [7:0] out1203;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1203 = in0;
    end

    reg [7:0] out1204;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1204 = in0;
    end

    reg [7:0] out1205;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1205 = in0;
    end

    reg [7:0] out1206;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1206 = in0;
    end

    reg [7:0] out1207;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1207 = in0;
    end

    reg [7:0] out1208;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1208 = in0;
    end

    reg [7:0] out1209;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1209 = in0;
    end

    reg [7:0] out1210;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1210 = in0;
    end

    reg [7:0] out1211;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1211 = in0;
    end

    reg [7:0] out1212;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1212 = in0;
    end

    reg [7:0] out1213;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1213 = in0;
    end

    reg [7:0] out1214;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1214 = in0;
    end

    reg [7:0] out1215;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1215 = in0;
    end

    reg [7:0] out1216;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1216 = in0;
    end

    reg [7:0] out1217;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1217 = in0;
    end

    reg [7:0] out1218;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1218 = in0;
    end

    reg [7:0] out1219;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1219 = in0;
    end

    reg [7:0] out1220;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1220 = in0;
    end

    reg [7:0] out1221;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1221 = in0;
    end

    reg [7:0] out1222;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1222 = in0;
    end

    reg [7:0] out1223;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1223 = in0;
    end

    reg [7:0] out1224;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1224 = in0;
    end

    reg [7:0] out1225;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1225 = in0;
    end

    reg [7:0] out1226;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1226 = in0;
    end

    reg [7:0] out1227;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1227 = in0;
    end

    reg [7:0] out1228;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1228 = in0;
    end

    reg [7:0] out1229;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1229 = in0;
    end

    reg [7:0] out1230;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1230 = in0;
    end

    reg [7:0] out1231;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1231 = in0;
    end

    reg [7:0] out1232;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1232 = in0;
    end

    reg [7:0] out1233;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1233 = in0;
    end

    reg [7:0] out1234;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1234 = in0;
    end

    reg [7:0] out1235;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1235 = in0;
    end

    reg [7:0] out1236;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1236 = in0;
    end

    reg [7:0] out1237;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1237 = in0;
    end

    reg [7:0] out1238;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1238 = in0;
    end

    reg [7:0] out1239;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1239 = in0;
    end

    reg [7:0] out1240;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1240 = in0;
    end

    reg [7:0] out1241;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1241 = in0;
    end

    reg [7:0] out1242;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1242 = in0;
    end

    reg [7:0] out1243;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1243 = in0;
    end

    reg [7:0] out1244;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1244 = in0;
    end

    reg [7:0] out1245;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1245 = in0;
    end

    reg [7:0] out1246;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1246 = in0;
    end

    reg [7:0] out1247;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1247 = in0;
    end

    reg [7:0] out1248;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1248 = in0;
    end

    reg [7:0] out1249;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1249 = in0;
    end

    reg [7:0] out1250;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1250 = in0;
    end

    reg [7:0] out1251;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1251 = in0;
    end

    reg [7:0] out1252;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1252 = in0;
    end

    reg [7:0] out1253;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1253 = in0;
    end

    reg [7:0] out1254;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1254 = in0;
    end

    reg [7:0] out1255;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1255 = in0;
    end

    reg [7:0] out1256;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1256 = in0;
    end

    reg [7:0] out1257;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1257 = in0;
    end

    reg [7:0] out1258;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1258 = in0;
    end

    reg [7:0] out1259;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1259 = in0;
    end

    reg [7:0] out1260;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1260 = in0;
    end

    reg [7:0] out1261;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1261 = in0;
    end

    reg [7:0] out1262;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1262 = in0;
    end

    reg [7:0] out1263;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1263 = in0;
    end

    reg [7:0] out1264;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1264 = in0;
    end

    reg [7:0] out1265;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1265 = in0;
    end

    reg [7:0] out1266;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1266 = in0;
    end

    reg [7:0] out1267;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1267 = in0;
    end

    reg [7:0] out1268;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1268 = in0;
    end

    reg [7:0] out1269;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1269 = in0;
    end

    reg [7:0] out1270;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1270 = in0;
    end

    reg [7:0] out1271;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1271 = in0;
    end

    reg [7:0] out1272;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1272 = in0;
    end

    reg [7:0] out1273;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1273 = in0;
    end

    reg [7:0] out1274;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1274 = in0;
    end

    reg [7:0] out1275;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1275 = in0;
    end

    reg [7:0] out1276;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1276 = in0;
    end

    reg [7:0] out1277;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1277 = in0;
    end

    reg [7:0] out1278;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1278 = in0;
    end

    reg [7:0] out1279;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1279 = in0;
    end

    reg [7:0] out1280;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1280 = in0;
    end

    reg [7:0] out1281;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1281 = in0;
    end

    reg [7:0] out1282;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1282 = in0;
    end

    reg [7:0] out1283;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1283 = in0;
    end

    reg [7:0] out1284;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1284 = in0;
    end

    reg [7:0] out1285;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1285 = in0;
    end

    reg [7:0] out1286;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1286 = in0;
    end

    reg [7:0] out1287;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1287 = in0;
    end

    reg [7:0] out1288;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1288 = in0;
    end

    reg [7:0] out1289;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1289 = in0;
    end

    reg [7:0] out1290;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1290 = in0;
    end

    reg [7:0] out1291;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1291 = in0;
    end

    reg [7:0] out1292;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1292 = in0;
    end

    reg [7:0] out1293;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1293 = in0;
    end

    reg [7:0] out1294;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1294 = in0;
    end

    reg [7:0] out1295;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1295 = in0;
    end

    reg [7:0] out1296;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1296 = in0;
    end

    reg [7:0] out1297;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1297 = in0;
    end

    reg [7:0] out1298;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1298 = in0;
    end

    reg [7:0] out1299;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1299 = in0;
    end

    reg [7:0] out1300;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1300 = in0;
    end

    reg [7:0] out1301;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1301 = in0;
    end

    reg [7:0] out1302;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1302 = in0;
    end

    reg [7:0] out1303;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1303 = in0;
    end

    reg [7:0] out1304;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1304 = in0;
    end

    reg [7:0] out1305;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1305 = in0;
    end

    reg [7:0] out1306;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1306 = in0;
    end

    reg [7:0] out1307;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1307 = in0;
    end

    reg [7:0] out1308;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1308 = in0;
    end

    reg [7:0] out1309;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1309 = in0;
    end

    reg [7:0] out1310;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1310 = in0;
    end

    reg [7:0] out1311;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1311 = in0;
    end

    reg [7:0] out1312;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1312 = in0;
    end

    reg [7:0] out1313;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1313 = in0;
    end

    reg [7:0] out1314;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1314 = in0;
    end

    reg [7:0] out1315;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1315 = in0;
    end

    reg [7:0] out1316;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1316 = in0;
    end

    reg [7:0] out1317;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1317 = in0;
    end

    reg [7:0] out1318;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1318 = in0;
    end

    reg [7:0] out1319;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1319 = in0;
    end

    reg [7:0] out1320;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1320 = in0;
    end

    reg [7:0] out1321;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1321 = in0;
    end

    reg [7:0] out1322;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1322 = in0;
    end

    reg [7:0] out1323;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1323 = in0;
    end

    reg [7:0] out1324;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1324 = in0;
    end

    reg [7:0] out1325;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1325 = in0;
    end

    reg [7:0] out1326;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1326 = in0;
    end

    reg [7:0] out1327;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1327 = in0;
    end

    reg [7:0] out1328;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1328 = in0;
    end

    reg [7:0] out1329;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1329 = in0;
    end

    reg [7:0] out1330;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1330 = in0;
    end

    reg [7:0] out1331;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1331 = in0;
    end

    reg [7:0] out1332;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1332 = in0;
    end

    reg [7:0] out1333;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1333 = in0;
    end

    reg [7:0] out1334;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1334 = in0;
    end

    reg [7:0] out1335;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1335 = in0;
    end

    reg [7:0] out1336;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1336 = in0;
    end

    reg [7:0] out1337;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1337 = in0;
    end

    reg [7:0] out1338;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1338 = in0;
    end

    reg [7:0] out1339;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1339 = in0;
    end

    reg [7:0] out1340;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1340 = in0;
    end

    reg [7:0] out1341;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1341 = in0;
    end

    reg [7:0] out1342;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1342 = in0;
    end

    reg [7:0] out1343;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1343 = in0;
    end

    reg [7:0] out1344;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1344 = in0;
    end

    reg [7:0] out1345;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1345 = in0;
    end

    reg [7:0] out1346;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1346 = in0;
    end

    reg [7:0] out1347;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1347 = in0;
    end

    reg [7:0] out1348;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1348 = in0;
    end

    reg [7:0] out1349;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1349 = in0;
    end

    reg [7:0] out1350;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1350 = in0;
    end

    reg [7:0] out1351;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1351 = in0;
    end

    reg [7:0] out1352;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1352 = in0;
    end

    reg [7:0] out1353;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1353 = in0;
    end

    reg [7:0] out1354;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1354 = in0;
    end

    reg [7:0] out1355;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1355 = in0;
    end

    reg [7:0] out1356;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1356 = in0;
    end

    reg [7:0] out1357;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1357 = in0;
    end

    reg [7:0] out1358;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1358 = in0;
    end

    reg [7:0] out1359;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1359 = in0;
    end

    reg [7:0] out1360;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1360 = in0;
    end

    reg [7:0] out1361;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1361 = in0;
    end

    reg [7:0] out1362;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1362 = in0;
    end

    reg [7:0] out1363;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1363 = in0;
    end

    reg [7:0] out1364;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1364 = in0;
    end

    reg [7:0] out1365;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1365 = in0;
    end

    reg [7:0] out1366;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1366 = in0;
    end

    reg [7:0] out1367;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1367 = in0;
    end

    reg [7:0] out1368;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1368 = in0;
    end

    reg [7:0] out1369;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1369 = in0;
    end

    reg [7:0] out1370;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1370 = in0;
    end

    reg [7:0] out1371;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1371 = in0;
    end

    reg [7:0] out1372;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1372 = in0;
    end

    reg [7:0] out1373;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1373 = in0;
    end

    reg [7:0] out1374;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1374 = in0;
    end

    reg [7:0] out1375;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1375 = in0;
    end

    reg [7:0] out1376;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1376 = in0;
    end

    reg [7:0] out1377;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1377 = in0;
    end

    reg [7:0] out1378;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1378 = in0;
    end

    reg [7:0] out1379;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1379 = in0;
    end

    reg [7:0] out1380;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1380 = in0;
    end

    reg [7:0] out1381;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1381 = in0;
    end

    reg [7:0] out1382;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1382 = in0;
    end

    reg [7:0] out1383;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1383 = in0;
    end

    reg [7:0] out1384;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1384 = in0;
    end

    reg [7:0] out1385;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1385 = in0;
    end

    reg [7:0] out1386;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1386 = in0;
    end

    reg [7:0] out1387;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1387 = in0;
    end

    reg [7:0] out1388;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1388 = in0;
    end

    reg [7:0] out1389;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1389 = in0;
    end

    reg [7:0] out1390;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1390 = in0;
    end

    reg [7:0] out1391;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1391 = in0;
    end

    reg [7:0] out1392;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1392 = in0;
    end

    reg [7:0] out1393;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1393 = in0;
    end

    reg [7:0] out1394;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1394 = in0;
    end

    reg [7:0] out1395;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1395 = in0;
    end

    reg [7:0] out1396;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1396 = in0;
    end

    reg [7:0] out1397;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1397 = in0;
    end

    reg [7:0] out1398;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1398 = in0;
    end

    reg [7:0] out1399;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1399 = in0;
    end

    reg [7:0] out1400;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1400 = in0;
    end

    reg [7:0] out1401;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1401 = in0;
    end

    reg [7:0] out1402;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1402 = in0;
    end

    reg [7:0] out1403;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1403 = in0;
    end

    reg [7:0] out1404;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1404 = in0;
    end

    reg [7:0] out1405;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1405 = in0;
    end

    reg [7:0] out1406;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1406 = in0;
    end

    reg [7:0] out1407;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1407 = in0;
    end

    reg [7:0] out1408;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1408 = in0;
    end

    reg [7:0] out1409;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1409 = in0;
    end

    reg [7:0] out1410;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1410 = in0;
    end

    reg [7:0] out1411;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1411 = in0;
    end

    reg [7:0] out1412;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1412 = in0;
    end

    reg [7:0] out1413;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1413 = in0;
    end

    reg [7:0] out1414;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1414 = in0;
    end

    reg [7:0] out1415;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1415 = in0;
    end

    reg [7:0] out1416;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1416 = in0;
    end

    reg [7:0] out1417;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1417 = in0;
    end

    reg [7:0] out1418;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1418 = in0;
    end

    reg [7:0] out1419;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1419 = in0;
    end

    reg [7:0] out1420;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1420 = in0;
    end

    reg [7:0] out1421;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1421 = in0;
    end

    reg [7:0] out1422;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1422 = in0;
    end

    reg [7:0] out1423;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1423 = in0;
    end

    reg [7:0] out1424;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1424 = in0;
    end

    reg [7:0] out1425;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1425 = in0;
    end

    reg [7:0] out1426;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1426 = in0;
    end

    reg [7:0] out1427;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1427 = in0;
    end

    reg [7:0] out1428;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1428 = in0;
    end

    reg [7:0] out1429;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1429 = in0;
    end

    reg [7:0] out1430;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1430 = in0;
    end

    reg [7:0] out1431;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1431 = in0;
    end

    reg [7:0] out1432;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1432 = in0;
    end

    reg [7:0] out1433;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1433 = in0;
    end

    reg [7:0] out1434;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1434 = in0;
    end

    reg [7:0] out1435;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1435 = in0;
    end

    reg [7:0] out1436;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1436 = in0;
    end

    reg [7:0] out1437;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1437 = in0;
    end

    reg [7:0] out1438;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1438 = in0;
    end

    reg [7:0] out1439;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1439 = in0;
    end

    reg [7:0] out1440;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1440 = in0;
    end

    reg [7:0] out1441;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1441 = in0;
    end

    reg [7:0] out1442;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1442 = in0;
    end

    reg [7:0] out1443;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1443 = in0;
    end

    reg [7:0] out1444;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1444 = in0;
    end

    reg [7:0] out1445;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1445 = in0;
    end

    reg [7:0] out1446;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1446 = in0;
    end

    reg [7:0] out1447;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1447 = in0;
    end

    reg [7:0] out1448;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1448 = in0;
    end

    reg [7:0] out1449;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1449 = in0;
    end

    reg [7:0] out1450;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1450 = in0;
    end

    reg [7:0] out1451;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1451 = in0;
    end

    reg [7:0] out1452;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1452 = in0;
    end

    reg [7:0] out1453;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1453 = in0;
    end

    reg [7:0] out1454;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1454 = in0;
    end

    reg [7:0] out1455;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1455 = in0;
    end

    reg [7:0] out1456;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1456 = in0;
    end

    reg [7:0] out1457;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1457 = in0;
    end

    reg [7:0] out1458;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1458 = in0;
    end

    reg [7:0] out1459;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1459 = in0;
    end

    reg [7:0] out1460;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1460 = in0;
    end

    reg [7:0] out1461;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1461 = in0;
    end

    reg [7:0] out1462;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1462 = in0;
    end

    reg [7:0] out1463;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1463 = in0;
    end

    reg [7:0] out1464;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1464 = in0;
    end

    reg [7:0] out1465;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1465 = in0;
    end

    reg [7:0] out1466;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1466 = in0;
    end

    reg [7:0] out1467;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1467 = in0;
    end

    reg [7:0] out1468;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1468 = in0;
    end

    reg [7:0] out1469;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1469 = in0;
    end

    reg [7:0] out1470;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1470 = in0;
    end

    reg [7:0] out1471;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1471 = in0;
    end

    reg [7:0] out1472;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1472 = in0;
    end

    reg [7:0] out1473;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1473 = in0;
    end

    reg [7:0] out1474;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1474 = in0;
    end

    reg [7:0] out1475;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1475 = in0;
    end

    reg [7:0] out1476;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1476 = in0;
    end

    reg [7:0] out1477;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1477 = in0;
    end

    reg [7:0] out1478;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1478 = in0;
    end

    reg [7:0] out1479;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1479 = in0;
    end

    reg [7:0] out1480;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1480 = in0;
    end

    reg [7:0] out1481;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1481 = in0;
    end

    reg [7:0] out1482;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1482 = in0;
    end

    reg [7:0] out1483;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1483 = in0;
    end

    reg [7:0] out1484;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1484 = in0;
    end

    reg [7:0] out1485;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1485 = in0;
    end

    reg [7:0] out1486;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1486 = in0;
    end

    reg [7:0] out1487;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1487 = in0;
    end

    reg [7:0] out1488;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1488 = in0;
    end

    reg [7:0] out1489;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1489 = in0;
    end

    reg [7:0] out1490;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1490 = in0;
    end

    reg [7:0] out1491;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1491 = in0;
    end

    reg [7:0] out1492;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1492 = in0;
    end

    reg [7:0] out1493;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1493 = in0;
    end

    reg [7:0] out1494;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1494 = in0;
    end

    reg [7:0] out1495;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1495 = in0;
    end

    reg [7:0] out1496;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1496 = in0;
    end

    reg [7:0] out1497;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1497 = in0;
    end

    reg [7:0] out1498;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1498 = in0;
    end

    reg [7:0] out1499;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1499 = in0;
    end

    reg [7:0] out1500;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1500 = in0;
    end

    reg [7:0] out1501;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1501 = in0;
    end

    reg [7:0] out1502;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1502 = in0;
    end

    reg [7:0] out1503;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1503 = in0;
    end

    reg [7:0] out1504;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1504 = in0;
    end

    reg [7:0] out1505;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1505 = in0;
    end

    reg [7:0] out1506;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1506 = in0;
    end

    reg [7:0] out1507;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1507 = in0;
    end

    reg [7:0] out1508;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1508 = in0;
    end

    reg [7:0] out1509;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1509 = in0;
    end

    reg [7:0] out1510;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1510 = in0;
    end

    reg [7:0] out1511;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1511 = in0;
    end

    reg [7:0] out1512;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1512 = in0;
    end

    reg [7:0] out1513;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1513 = in0;
    end

    reg [7:0] out1514;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1514 = in0;
    end

    reg [7:0] out1515;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1515 = in0;
    end

    reg [7:0] out1516;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1516 = in0;
    end

    reg [7:0] out1517;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1517 = in0;
    end

    reg [7:0] out1518;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1518 = in0;
    end

    reg [7:0] out1519;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1519 = in0;
    end

    reg [7:0] out1520;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1520 = in0;
    end

    reg [7:0] out1521;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1521 = in0;
    end

    reg [7:0] out1522;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1522 = in0;
    end

    reg [7:0] out1523;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1523 = in0;
    end

    reg [7:0] out1524;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1524 = in0;
    end

    reg [7:0] out1525;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1525 = in0;
    end

    reg [7:0] out1526;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1526 = in0;
    end

    reg [7:0] out1527;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1527 = in0;
    end

    reg [7:0] out1528;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1528 = in0;
    end

    reg [7:0] out1529;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1529 = in0;
    end

    reg [7:0] out1530;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1530 = in0;
    end

    reg [7:0] out1531;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1531 = in0;
    end

    reg [7:0] out1532;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1532 = in0;
    end

    reg [7:0] out1533;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1533 = in0;
    end

    reg [7:0] out1534;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1534 = in0;
    end

    reg [7:0] out1535;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1535 = in0;
    end

    reg [7:0] out1536;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1536 = in0;
    end

    reg [7:0] out1537;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1537 = in0;
    end

    reg [7:0] out1538;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1538 = in0;
    end

    reg [7:0] out1539;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1539 = in0;
    end

    reg [7:0] out1540;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1540 = in0;
    end

    reg [7:0] out1541;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1541 = in0;
    end

    reg [7:0] out1542;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1542 = in0;
    end

    reg [7:0] out1543;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1543 = in0;
    end

    reg [7:0] out1544;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1544 = in0;
    end

    reg [7:0] out1545;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1545 = in0;
    end

    reg [7:0] out1546;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1546 = in0;
    end

    reg [7:0] out1547;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1547 = in0;
    end

    reg [7:0] out1548;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1548 = in0;
    end

    reg [7:0] out1549;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1549 = in0;
    end

    reg [7:0] out1550;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1550 = in0;
    end

    reg [7:0] out1551;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1551 = in0;
    end

    reg [7:0] out1552;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1552 = in0;
    end

    reg [7:0] out1553;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1553 = in0;
    end

    reg [7:0] out1554;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1554 = in0;
    end

    reg [7:0] out1555;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1555 = in0;
    end

    reg [7:0] out1556;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1556 = in0;
    end

    reg [7:0] out1557;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1557 = in0;
    end

    reg [7:0] out1558;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1558 = in0;
    end

    reg [7:0] out1559;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1559 = in0;
    end

    reg [7:0] out1560;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1560 = in0;
    end

    reg [7:0] out1561;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1561 = in0;
    end

    reg [7:0] out1562;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1562 = in0;
    end

    reg [7:0] out1563;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1563 = in0;
    end

    reg [7:0] out1564;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1564 = in0;
    end

    reg [7:0] out1565;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1565 = in0;
    end

    reg [7:0] out1566;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1566 = in0;
    end

    reg [7:0] out1567;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1567 = in0;
    end

    reg [7:0] out1568;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1568 = in0;
    end

    reg [7:0] out1569;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1569 = in0;
    end

    reg [7:0] out1570;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1570 = in0;
    end

    reg [7:0] out1571;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1571 = in0;
    end

    reg [7:0] out1572;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1572 = in0;
    end

    reg [7:0] out1573;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1573 = in0;
    end

    reg [7:0] out1574;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1574 = in0;
    end

    reg [7:0] out1575;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1575 = in0;
    end

    reg [7:0] out1576;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1576 = in0;
    end

    reg [7:0] out1577;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1577 = in0;
    end

    reg [7:0] out1578;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1578 = in0;
    end

    reg [7:0] out1579;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1579 = in0;
    end

    reg [7:0] out1580;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1580 = in0;
    end

    reg [7:0] out1581;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1581 = in0;
    end

    reg [7:0] out1582;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1582 = in0;
    end

    reg [7:0] out1583;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1583 = in0;
    end

    reg [7:0] out1584;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1584 = in0;
    end

    reg [7:0] out1585;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1585 = in0;
    end

    reg [7:0] out1586;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1586 = in0;
    end

    reg [7:0] out1587;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1587 = in0;
    end

    reg [7:0] out1588;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1588 = in0;
    end

    reg [7:0] out1589;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1589 = in0;
    end

    reg [7:0] out1590;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1590 = in0;
    end

    reg [7:0] out1591;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1591 = in0;
    end

    reg [7:0] out1592;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1592 = in0;
    end

    reg [7:0] out1593;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1593 = in0;
    end

    reg [7:0] out1594;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1594 = in0;
    end

    reg [7:0] out1595;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1595 = in0;
    end

    reg [7:0] out1596;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1596 = in0;
    end

    reg [7:0] out1597;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1597 = in0;
    end

    reg [7:0] out1598;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1598 = in0;
    end

    reg [7:0] out1599;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1599 = in0;
    end

    reg [7:0] out1600;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1600 = in0;
    end

    reg [7:0] out1601;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1601 = in0;
    end

    reg [7:0] out1602;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1602 = in0;
    end

    reg [7:0] out1603;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1603 = in0;
    end

    reg [7:0] out1604;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1604 = in0;
    end

    reg [7:0] out1605;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1605 = in0;
    end

    reg [7:0] out1606;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1606 = in0;
    end

    reg [7:0] out1607;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1607 = in0;
    end

    reg [7:0] out1608;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1608 = in0;
    end

    reg [7:0] out1609;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1609 = in0;
    end

    reg [7:0] out1610;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1610 = in0;
    end

    reg [7:0] out1611;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1611 = in0;
    end

    reg [7:0] out1612;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1612 = in0;
    end

    reg [7:0] out1613;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1613 = in0;
    end

    reg [7:0] out1614;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1614 = in0;
    end

    reg [7:0] out1615;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1615 = in0;
    end

    reg [7:0] out1616;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1616 = in0;
    end

    reg [7:0] out1617;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1617 = in0;
    end

    reg [7:0] out1618;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1618 = in0;
    end

    reg [7:0] out1619;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1619 = in0;
    end

    reg [7:0] out1620;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1620 = in0;
    end

    reg [7:0] out1621;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1621 = in0;
    end

    reg [7:0] out1622;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1622 = in0;
    end

    reg [7:0] out1623;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1623 = in0;
    end

    reg [7:0] out1624;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1624 = in0;
    end

    reg [7:0] out1625;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1625 = in0;
    end

    reg [7:0] out1626;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1626 = in0;
    end

    reg [7:0] out1627;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1627 = in0;
    end

    reg [7:0] out1628;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1628 = in0;
    end

    reg [7:0] out1629;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1629 = in0;
    end

    reg [7:0] out1630;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1630 = in0;
    end

    reg [7:0] out1631;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1631 = in0;
    end

    reg [7:0] out1632;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1632 = in0;
    end

    reg [7:0] out1633;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1633 = in0;
    end

    reg [7:0] out1634;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1634 = in0;
    end

    reg [7:0] out1635;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1635 = in0;
    end

    reg [7:0] out1636;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1636 = in0;
    end

    reg [7:0] out1637;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1637 = in0;
    end

    reg [7:0] out1638;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1638 = in0;
    end

    reg [7:0] out1639;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1639 = in0;
    end

    reg [7:0] out1640;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1640 = in0;
    end

    reg [7:0] out1641;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1641 = in0;
    end

    reg [7:0] out1642;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1642 = in0;
    end

    reg [7:0] out1643;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1643 = in0;
    end

    reg [7:0] out1644;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1644 = in0;
    end

    reg [7:0] out1645;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1645 = in0;
    end

    reg [7:0] out1646;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1646 = in0;
    end

    reg [7:0] out1647;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1647 = in0;
    end

    reg [7:0] out1648;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1648 = in0;
    end

    reg [7:0] out1649;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1649 = in0;
    end

    reg [7:0] out1650;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1650 = in0;
    end

    reg [7:0] out1651;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1651 = in0;
    end

    reg [7:0] out1652;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1652 = in0;
    end

    reg [7:0] out1653;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1653 = in0;
    end

    reg [7:0] out1654;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1654 = in0;
    end

    reg [7:0] out1655;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1655 = in0;
    end

    reg [7:0] out1656;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1656 = in0;
    end

    reg [7:0] out1657;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1657 = in0;
    end

    reg [7:0] out1658;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1658 = in0;
    end

    reg [7:0] out1659;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1659 = in0;
    end

    reg [7:0] out1660;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1660 = in0;
    end

    reg [7:0] out1661;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1661 = in0;
    end

    reg [7:0] out1662;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1662 = in0;
    end

    reg [7:0] out1663;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1663 = in0;
    end

    reg [7:0] out1664;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1664 = in0;
    end

    reg [7:0] out1665;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1665 = in0;
    end

    reg [7:0] out1666;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1666 = in0;
    end

    reg [7:0] out1667;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1667 = in0;
    end

    reg [7:0] out1668;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1668 = in0;
    end

    reg [7:0] out1669;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1669 = in0;
    end

    reg [7:0] out1670;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1670 = in0;
    end

    reg [7:0] out1671;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1671 = in0;
    end

    reg [7:0] out1672;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1672 = in0;
    end

    reg [7:0] out1673;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1673 = in0;
    end

    reg [7:0] out1674;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1674 = in0;
    end

    reg [7:0] out1675;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1675 = in0;
    end

    reg [7:0] out1676;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1676 = in0;
    end

    reg [7:0] out1677;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1677 = in0;
    end

    reg [7:0] out1678;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1678 = in0;
    end

    reg [7:0] out1679;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1679 = in0;
    end

    reg [7:0] out1680;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1680 = in0;
    end

    reg [7:0] out1681;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1681 = in0;
    end

    reg [7:0] out1682;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1682 = in0;
    end

    reg [7:0] out1683;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1683 = in0;
    end

    reg [7:0] out1684;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1684 = in0;
    end

    reg [7:0] out1685;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1685 = in0;
    end

    reg [7:0] out1686;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1686 = in0;
    end

    reg [7:0] out1687;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1687 = in0;
    end

    reg [7:0] out1688;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1688 = in0;
    end

    reg [7:0] out1689;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1689 = in0;
    end

    reg [7:0] out1690;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1690 = in0;
    end

    reg [7:0] out1691;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1691 = in0;
    end

    reg [7:0] out1692;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1692 = in0;
    end

    reg [7:0] out1693;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1693 = in0;
    end

    reg [7:0] out1694;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1694 = in0;
    end

    reg [7:0] out1695;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1695 = in0;
    end

    reg [7:0] out1696;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1696 = in0;
    end

    reg [7:0] out1697;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1697 = in0;
    end

    reg [7:0] out1698;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1698 = in0;
    end

    reg [7:0] out1699;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1699 = in0;
    end

    reg [7:0] out1700;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1700 = in0;
    end

    reg [7:0] out1701;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1701 = in0;
    end

    reg [7:0] out1702;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1702 = in0;
    end

    reg [7:0] out1703;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1703 = in0;
    end

    reg [7:0] out1704;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1704 = in0;
    end

    reg [7:0] out1705;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1705 = in0;
    end

    reg [7:0] out1706;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1706 = in0;
    end

    reg [7:0] out1707;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1707 = in0;
    end

    reg [7:0] out1708;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1708 = in0;
    end

    reg [7:0] out1709;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1709 = in0;
    end

    reg [7:0] out1710;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1710 = in0;
    end

    reg [7:0] out1711;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1711 = in0;
    end

    reg [7:0] out1712;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1712 = in0;
    end

    reg [7:0] out1713;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1713 = in0;
    end

    reg [7:0] out1714;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1714 = in0;
    end

    reg [7:0] out1715;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1715 = in0;
    end

    reg [7:0] out1716;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1716 = in0;
    end

    reg [7:0] out1717;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1717 = in0;
    end

    reg [7:0] out1718;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1718 = in0;
    end

    reg [7:0] out1719;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1719 = in0;
    end

    reg [7:0] out1720;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1720 = in0;
    end

    reg [7:0] out1721;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1721 = in0;
    end

    reg [7:0] out1722;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1722 = in0;
    end

    reg [7:0] out1723;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1723 = in0;
    end

    reg [7:0] out1724;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1724 = in0;
    end

    reg [7:0] out1725;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1725 = in0;
    end

    reg [7:0] out1726;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1726 = in0;
    end

    reg [7:0] out1727;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1727 = in0;
    end

    reg [7:0] out1728;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1728 = in0;
    end

    reg [7:0] out1729;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1729 = in0;
    end

    reg [7:0] out1730;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1730 = in0;
    end

    reg [7:0] out1731;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1731 = in0;
    end

    reg [7:0] out1732;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1732 = in0;
    end

    reg [7:0] out1733;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1733 = in0;
    end

    reg [7:0] out1734;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1734 = in0;
    end

    reg [7:0] out1735;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1735 = in0;
    end

    reg [7:0] out1736;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1736 = in0;
    end

    reg [7:0] out1737;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1737 = in0;
    end

    reg [7:0] out1738;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1738 = in0;
    end

    reg [7:0] out1739;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1739 = in0;
    end

    reg [7:0] out1740;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1740 = in0;
    end

    reg [7:0] out1741;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1741 = in0;
    end

    reg [7:0] out1742;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1742 = in0;
    end

    reg [7:0] out1743;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1743 = in0;
    end

    reg [7:0] out1744;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1744 = in0;
    end

    reg [7:0] out1745;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1745 = in0;
    end

    reg [7:0] out1746;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1746 = in0;
    end

    reg [7:0] out1747;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1747 = in0;
    end

    reg [7:0] out1748;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1748 = in0;
    end

    reg [7:0] out1749;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1749 = in0;
    end

    reg [7:0] out1750;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1750 = in0;
    end

    reg [7:0] out1751;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1751 = in0;
    end

    reg [7:0] out1752;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1752 = in0;
    end

    reg [7:0] out1753;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1753 = in0;
    end

    reg [7:0] out1754;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1754 = in0;
    end

    reg [7:0] out1755;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1755 = in0;
    end

    reg [7:0] out1756;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1756 = in0;
    end

    reg [7:0] out1757;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1757 = in0;
    end

    reg [7:0] out1758;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1758 = in0;
    end

    reg [7:0] out1759;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1759 = in0;
    end

    reg [7:0] out1760;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1760 = in0;
    end

    reg [7:0] out1761;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1761 = in0;
    end

    reg [7:0] out1762;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1762 = in0;
    end

    reg [7:0] out1763;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1763 = in0;
    end

    reg [7:0] out1764;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1764 = in0;
    end

    reg [7:0] out1765;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1765 = in0;
    end

    reg [7:0] out1766;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1766 = in0;
    end

    reg [7:0] out1767;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1767 = in0;
    end

    reg [7:0] out1768;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1768 = in0;
    end

    reg [7:0] out1769;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1769 = in0;
    end

    reg [7:0] out1770;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1770 = in0;
    end

    reg [7:0] out1771;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1771 = in0;
    end

    reg [7:0] out1772;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1772 = in0;
    end

    reg [7:0] out1773;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1773 = in0;
    end

    reg [7:0] out1774;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1774 = in0;
    end

    reg [7:0] out1775;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1775 = in0;
    end

    reg [7:0] out1776;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1776 = in0;
    end

    reg [7:0] out1777;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1777 = in0;
    end

    reg [7:0] out1778;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1778 = in0;
    end

    reg [7:0] out1779;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1779 = in0;
    end

    reg [7:0] out1780;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1780 = in0;
    end

    reg [7:0] out1781;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1781 = in0;
    end

    reg [7:0] out1782;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1782 = in0;
    end

    reg [7:0] out1783;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1783 = in0;
    end

    reg [7:0] out1784;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1784 = in0;
    end

    reg [7:0] out1785;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1785 = in0;
    end

    reg [7:0] out1786;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1786 = in0;
    end

    reg [7:0] out1787;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1787 = in0;
    end

    reg [7:0] out1788;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1788 = in0;
    end

    reg [7:0] out1789;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1789 = in0;
    end

    reg [7:0] out1790;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1790 = in0;
    end

    reg [7:0] out1791;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1791 = in0;
    end

    reg [7:0] out1792;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1792 = in0;
    end

    reg [7:0] out1793;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1793 = in0;
    end

    reg [7:0] out1794;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1794 = in0;
    end

    reg [7:0] out1795;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1795 = in0;
    end

    reg [7:0] out1796;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1796 = in0;
    end

    reg [7:0] out1797;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1797 = in0;
    end

    reg [7:0] out1798;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1798 = in0;
    end

    reg [7:0] out1799;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1799 = in0;
    end

    reg [7:0] out1800;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1800 = in0;
    end

    reg [7:0] out1801;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1801 = in0;
    end

    reg [7:0] out1802;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1802 = in0;
    end

    reg [7:0] out1803;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1803 = in0;
    end

    reg [7:0] out1804;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1804 = in0;
    end

    reg [7:0] out1805;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1805 = in0;
    end

    reg [7:0] out1806;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1806 = in0;
    end

    reg [7:0] out1807;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1807 = in0;
    end

    reg [7:0] out1808;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1808 = in0;
    end

    reg [7:0] out1809;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1809 = in0;
    end

    reg [7:0] out1810;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1810 = in0;
    end

    reg [7:0] out1811;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1811 = in0;
    end

    reg [7:0] out1812;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1812 = in0;
    end

    reg [7:0] out1813;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1813 = in0;
    end

    reg [7:0] out1814;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1814 = in0;
    end

    reg [7:0] out1815;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1815 = in0;
    end

    reg [7:0] out1816;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1816 = in0;
    end

    reg [7:0] out1817;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1817 = in0;
    end

    reg [7:0] out1818;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1818 = in0;
    end

    reg [7:0] out1819;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1819 = in0;
    end

    reg [7:0] out1820;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1820 = in0;
    end

    reg [7:0] out1821;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1821 = in0;
    end

    reg [7:0] out1822;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1822 = in0;
    end

    reg [7:0] out1823;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1823 = in0;
    end

    reg [7:0] out1824;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1824 = in0;
    end

    reg [7:0] out1825;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1825 = in0;
    end

    reg [7:0] out1826;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1826 = in0;
    end

    reg [7:0] out1827;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1827 = in0;
    end

    reg [7:0] out1828;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1828 = in0;
    end

    reg [7:0] out1829;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1829 = in0;
    end

    reg [7:0] out1830;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1830 = in0;
    end

    reg [7:0] out1831;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1831 = in0;
    end

    reg [7:0] out1832;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1832 = in0;
    end

    reg [7:0] out1833;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1833 = in0;
    end

    reg [7:0] out1834;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1834 = in0;
    end

    reg [7:0] out1835;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1835 = in0;
    end

    reg [7:0] out1836;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1836 = in0;
    end

    reg [7:0] out1837;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1837 = in0;
    end

    reg [7:0] out1838;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1838 = in0;
    end

    reg [7:0] out1839;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1839 = in0;
    end

    reg [7:0] out1840;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1840 = in0;
    end

    reg [7:0] out1841;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1841 = in0;
    end

    reg [7:0] out1842;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1842 = in0;
    end

    reg [7:0] out1843;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1843 = in0;
    end

    reg [7:0] out1844;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1844 = in0;
    end

    reg [7:0] out1845;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1845 = in0;
    end

    reg [7:0] out1846;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1846 = in0;
    end

    reg [7:0] out1847;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1847 = in0;
    end

    reg [7:0] out1848;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1848 = in0;
    end

    reg [7:0] out1849;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1849 = in0;
    end

    reg [7:0] out1850;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1850 = in0;
    end

    reg [7:0] out1851;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1851 = in0;
    end

    reg [7:0] out1852;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1852 = in0;
    end

    reg [7:0] out1853;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1853 = in0;
    end

    reg [7:0] out1854;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1854 = in0;
    end

    reg [7:0] out1855;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1855 = in0;
    end

    reg [7:0] out1856;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1856 = in0;
    end

    reg [7:0] out1857;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1857 = in0;
    end

    reg [7:0] out1858;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1858 = in0;
    end

    reg [7:0] out1859;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1859 = in0;
    end

    reg [7:0] out1860;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1860 = in0;
    end

    reg [7:0] out1861;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1861 = in0;
    end

    reg [7:0] out1862;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1862 = in0;
    end

    reg [7:0] out1863;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1863 = in0;
    end

    reg [7:0] out1864;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1864 = in0;
    end

    reg [7:0] out1865;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1865 = in0;
    end

    reg [7:0] out1866;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1866 = in0;
    end

    reg [7:0] out1867;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1867 = in0;
    end

    reg [7:0] out1868;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1868 = in0;
    end

    reg [7:0] out1869;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1869 = in0;
    end

    reg [7:0] out1870;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1870 = in0;
    end

    reg [7:0] out1871;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1871 = in0;
    end

    reg [7:0] out1872;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1872 = in0;
    end

    reg [7:0] out1873;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1873 = in0;
    end

    reg [7:0] out1874;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1874 = in0;
    end

    reg [7:0] out1875;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1875 = in0;
    end

    reg [7:0] out1876;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1876 = in0;
    end

    reg [7:0] out1877;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1877 = in0;
    end

    reg [7:0] out1878;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1878 = in0;
    end

    reg [7:0] out1879;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1879 = in0;
    end

    reg [7:0] out1880;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1880 = in0;
    end

    reg [7:0] out1881;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1881 = in0;
    end

    reg [7:0] out1882;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1882 = in0;
    end

    reg [7:0] out1883;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1883 = in0;
    end

    reg [7:0] out1884;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1884 = in0;
    end

    reg [7:0] out1885;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1885 = in0;
    end

    reg [7:0] out1886;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1886 = in0;
    end

    reg [7:0] out1887;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1887 = in0;
    end

    reg [7:0] out1888;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1888 = in0;
    end

    reg [7:0] out1889;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1889 = in0;
    end

    reg [7:0] out1890;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1890 = in0;
    end

    reg [7:0] out1891;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1891 = in0;
    end

    reg [7:0] out1892;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1892 = in0;
    end

    reg [7:0] out1893;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1893 = in0;
    end

    reg [7:0] out1894;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1894 = in0;
    end

    reg [7:0] out1895;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1895 = in0;
    end

    reg [7:0] out1896;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1896 = in0;
    end

    reg [7:0] out1897;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1897 = in0;
    end

    reg [7:0] out1898;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1898 = in0;
    end

    reg [7:0] out1899;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1899 = in0;
    end

    reg [7:0] out1900;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1900 = in0;
    end

    reg [7:0] out1901;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1901 = in0;
    end

    reg [7:0] out1902;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1902 = in0;
    end

    reg [7:0] out1903;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1903 = in0;
    end

    reg [7:0] out1904;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1904 = in0;
    end

    reg [7:0] out1905;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1905 = in0;
    end

    reg [7:0] out1906;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1906 = in0;
    end

    reg [7:0] out1907;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1907 = in0;
    end

    reg [7:0] out1908;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1908 = in0;
    end

    reg [7:0] out1909;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1909 = in0;
    end

    reg [7:0] out1910;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1910 = in0;
    end

    reg [7:0] out1911;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1911 = in0;
    end

    reg [7:0] out1912;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1912 = in0;
    end

    reg [7:0] out1913;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1913 = in0;
    end

    reg [7:0] out1914;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1914 = in0;
    end

    reg [7:0] out1915;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1915 = in0;
    end

    reg [7:0] out1916;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1916 = in0;
    end

    reg [7:0] out1917;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1917 = in0;
    end

    reg [7:0] out1918;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1918 = in0;
    end

    reg [7:0] out1919;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1919 = in0;
    end

    reg [7:0] out1920;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1920 = in0;
    end

    reg [7:0] out1921;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1921 = in0;
    end

    reg [7:0] out1922;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1922 = in0;
    end

    reg [7:0] out1923;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1923 = in0;
    end

    reg [7:0] out1924;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1924 = in0;
    end

    reg [7:0] out1925;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1925 = in0;
    end

    reg [7:0] out1926;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1926 = in0;
    end

    reg [7:0] out1927;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1927 = in0;
    end

    reg [7:0] out1928;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1928 = in0;
    end

    reg [7:0] out1929;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1929 = in0;
    end

    reg [7:0] out1930;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1930 = in0;
    end

    reg [7:0] out1931;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1931 = in0;
    end

    reg [7:0] out1932;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1932 = in0;
    end

    reg [7:0] out1933;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1933 = in0;
    end

    reg [7:0] out1934;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1934 = in0;
    end

    reg [7:0] out1935;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1935 = in0;
    end

    reg [7:0] out1936;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1936 = in0;
    end

    reg [7:0] out1937;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1937 = in0;
    end

    reg [7:0] out1938;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1938 = in0;
    end

    reg [7:0] out1939;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1939 = in0;
    end

    reg [7:0] out1940;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1940 = in0;
    end

    reg [7:0] out1941;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1941 = in0;
    end

    reg [7:0] out1942;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1942 = in0;
    end

    reg [7:0] out1943;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1943 = in0;
    end

    reg [7:0] out1944;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1944 = in0;
    end

    reg [7:0] out1945;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1945 = in0;
    end

    reg [7:0] out1946;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1946 = in0;
    end

    reg [7:0] out1947;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1947 = in0;
    end

    reg [7:0] out1948;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1948 = in0;
    end

    reg [7:0] out1949;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1949 = in0;
    end

    reg [7:0] out1950;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1950 = in0;
    end

    reg [7:0] out1951;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1951 = in0;
    end

    reg [7:0] out1952;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1952 = in0;
    end

    reg [7:0] out1953;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1953 = in0;
    end

    reg [7:0] out1954;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1954 = in0;
    end

    reg [7:0] out1955;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1955 = in0;
    end

    reg [7:0] out1956;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1956 = in0;
    end

    reg [7:0] out1957;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1957 = in0;
    end

    reg [7:0] out1958;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1958 = in0;
    end

    reg [7:0] out1959;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1959 = in0;
    end

    reg [7:0] out1960;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1960 = in0;
    end

    reg [7:0] out1961;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1961 = in0;
    end

    reg [7:0] out1962;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1962 = in0;
    end

    reg [7:0] out1963;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1963 = in0;
    end

    reg [7:0] out1964;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1964 = in0;
    end

    reg [7:0] out1965;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1965 = in0;
    end

    reg [7:0] out1966;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1966 = in0;
    end

    reg [7:0] out1967;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1967 = in0;
    end

    reg [7:0] out1968;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1968 = in0;
    end

    reg [7:0] out1969;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1969 = in0;
    end

    reg [7:0] out1970;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1970 = in0;
    end

    reg [7:0] out1971;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1971 = in0;
    end

    reg [7:0] out1972;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1972 = in0;
    end

    reg [7:0] out1973;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1973 = in0;
    end

    reg [7:0] out1974;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1974 = in0;
    end

    reg [7:0] out1975;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1975 = in0;
    end

    reg [7:0] out1976;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1976 = in0;
    end

    reg [7:0] out1977;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1977 = in0;
    end

    reg [7:0] out1978;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1978 = in0;
    end

    reg [7:0] out1979;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1979 = in0;
    end

    reg [7:0] out1980;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1980 = in0;
    end

    reg [7:0] out1981;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1981 = in0;
    end

    reg [7:0] out1982;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1982 = in0;
    end

    reg [7:0] out1983;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1983 = in0;
    end

    reg [7:0] out1984;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1984 = in0;
    end

    reg [7:0] out1985;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1985 = in0;
    end

    reg [7:0] out1986;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1986 = in0;
    end

    reg [7:0] out1987;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1987 = in0;
    end

    reg [7:0] out1988;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1988 = in0;
    end

    reg [7:0] out1989;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1989 = in0;
    end

    reg [7:0] out1990;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1990 = in0;
    end

    reg [7:0] out1991;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1991 = in0;
    end

    reg [7:0] out1992;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1992 = in0;
    end

    reg [7:0] out1993;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1993 = in0;
    end

    reg [7:0] out1994;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1994 = in0;
    end

    reg [7:0] out1995;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1995 = in0;
    end

    reg [7:0] out1996;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1996 = in0;
    end

    reg [7:0] out1997;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1997 = in0;
    end

    reg [7:0] out1998;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1998 = in0;
    end

    reg [7:0] out1999;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out1999 = in0;
    end

    reg [7:0] out2000;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2000 = in0;
    end

    reg [7:0] out2001;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2001 = in0;
    end

    reg [7:0] out2002;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2002 = in0;
    end

    reg [7:0] out2003;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2003 = in0;
    end

    reg [7:0] out2004;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2004 = in0;
    end

    reg [7:0] out2005;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2005 = in0;
    end

    reg [7:0] out2006;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2006 = in0;
    end

    reg [7:0] out2007;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2007 = in0;
    end

    reg [7:0] out2008;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2008 = in0;
    end

    reg [7:0] out2009;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2009 = in0;
    end

    reg [7:0] out2010;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2010 = in0;
    end

    reg [7:0] out2011;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2011 = in0;
    end

    reg [7:0] out2012;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2012 = in0;
    end

    reg [7:0] out2013;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2013 = in0;
    end

    reg [7:0] out2014;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2014 = in0;
    end

    reg [7:0] out2015;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2015 = in0;
    end

    reg [7:0] out2016;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2016 = in0;
    end

    reg [7:0] out2017;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2017 = in0;
    end

    reg [7:0] out2018;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2018 = in0;
    end

    reg [7:0] out2019;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2019 = in0;
    end

    reg [7:0] out2020;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2020 = in0;
    end

    reg [7:0] out2021;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2021 = in0;
    end

    reg [7:0] out2022;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2022 = in0;
    end

    reg [7:0] out2023;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2023 = in0;
    end

    reg [7:0] out2024;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2024 = in0;
    end

    reg [7:0] out2025;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2025 = in0;
    end

    reg [7:0] out2026;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2026 = in0;
    end

    reg [7:0] out2027;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2027 = in0;
    end

    reg [7:0] out2028;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2028 = in0;
    end

    reg [7:0] out2029;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2029 = in0;
    end

    reg [7:0] out2030;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2030 = in0;
    end

    reg [7:0] out2031;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2031 = in0;
    end

    reg [7:0] out2032;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2032 = in0;
    end

    reg [7:0] out2033;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2033 = in0;
    end

    reg [7:0] out2034;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2034 = in0;
    end

    reg [7:0] out2035;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2035 = in0;
    end

    reg [7:0] out2036;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2036 = in0;
    end

    reg [7:0] out2037;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2037 = in0;
    end

    reg [7:0] out2038;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2038 = in0;
    end

    reg [7:0] out2039;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2039 = in0;
    end

    reg [7:0] out2040;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2040 = in0;
    end

    reg [7:0] out2041;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2041 = in0;
    end

    reg [7:0] out2042;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2042 = in0;
    end

    reg [7:0] out2043;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2043 = in0;
    end

    reg [7:0] out2044;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2044 = in0;
    end

    reg [7:0] out2045;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2045 = in0;
    end

    reg [7:0] out2046;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2046 = in0;
    end

    reg [7:0] out2047;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2047 = in0;
    end

    reg [7:0] out2048;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2048 = in0;
    end

    reg [7:0] out2049;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2049 = in0;
    end

    reg [7:0] out2050;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2050 = in0;
    end

    reg [7:0] out2051;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2051 = in0;
    end

    reg [7:0] out2052;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2052 = in0;
    end

    reg [7:0] out2053;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2053 = in0;
    end

    reg [7:0] out2054;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2054 = in0;
    end

    reg [7:0] out2055;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2055 = in0;
    end

    reg [7:0] out2056;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2056 = in0;
    end

    reg [7:0] out2057;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2057 = in0;
    end

    reg [7:0] out2058;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2058 = in0;
    end

    reg [7:0] out2059;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2059 = in0;
    end

    reg [7:0] out2060;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2060 = in0;
    end

    reg [7:0] out2061;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2061 = in0;
    end

    reg [7:0] out2062;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2062 = in0;
    end

    reg [7:0] out2063;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2063 = in0;
    end

    reg [7:0] out2064;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2064 = in0;
    end

    reg [7:0] out2065;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2065 = in0;
    end

    reg [7:0] out2066;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2066 = in0;
    end

    reg [7:0] out2067;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2067 = in0;
    end

    reg [7:0] out2068;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2068 = in0;
    end

    reg [7:0] out2069;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2069 = in0;
    end

    reg [7:0] out2070;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2070 = in0;
    end

    reg [7:0] out2071;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2071 = in0;
    end

    reg [7:0] out2072;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2072 = in0;
    end

    reg [7:0] out2073;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2073 = in0;
    end

    reg [7:0] out2074;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2074 = in0;
    end

    reg [7:0] out2075;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2075 = in0;
    end

    reg [7:0] out2076;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2076 = in0;
    end

    reg [7:0] out2077;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2077 = in0;
    end

    reg [7:0] out2078;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2078 = in0;
    end

    reg [7:0] out2079;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2079 = in0;
    end

    reg [7:0] out2080;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2080 = in0;
    end

    reg [7:0] out2081;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2081 = in0;
    end

    reg [7:0] out2082;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2082 = in0;
    end

    reg [7:0] out2083;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2083 = in0;
    end

    reg [7:0] out2084;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2084 = in0;
    end

    reg [7:0] out2085;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2085 = in0;
    end

    reg [7:0] out2086;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2086 = in0;
    end

    reg [7:0] out2087;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2087 = in0;
    end

    reg [7:0] out2088;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2088 = in0;
    end

    reg [7:0] out2089;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2089 = in0;
    end

    reg [7:0] out2090;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2090 = in0;
    end

    reg [7:0] out2091;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2091 = in0;
    end

    reg [7:0] out2092;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2092 = in0;
    end

    reg [7:0] out2093;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2093 = in0;
    end

    reg [7:0] out2094;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2094 = in0;
    end

    reg [7:0] out2095;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2095 = in0;
    end

    reg [7:0] out2096;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2096 = in0;
    end

    reg [7:0] out2097;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2097 = in0;
    end

    reg [7:0] out2098;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2098 = in0;
    end

    reg [7:0] out2099;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2099 = in0;
    end

    reg [7:0] out2100;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2100 = in0;
    end

    reg [7:0] out2101;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2101 = in0;
    end

    reg [7:0] out2102;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2102 = in0;
    end

    reg [7:0] out2103;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2103 = in0;
    end

    reg [7:0] out2104;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2104 = in0;
    end

    reg [7:0] out2105;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2105 = in0;
    end

    reg [7:0] out2106;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2106 = in0;
    end

    reg [7:0] out2107;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2107 = in0;
    end

    reg [7:0] out2108;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2108 = in0;
    end

    reg [7:0] out2109;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2109 = in0;
    end

    reg [7:0] out2110;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2110 = in0;
    end

    reg [7:0] out2111;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2111 = in0;
    end

    reg [7:0] out2112;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2112 = in0;
    end

    reg [7:0] out2113;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2113 = in0;
    end

    reg [7:0] out2114;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2114 = in0;
    end

    reg [7:0] out2115;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2115 = in0;
    end

    reg [7:0] out2116;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2116 = in0;
    end

    reg [7:0] out2117;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2117 = in0;
    end

    reg [7:0] out2118;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2118 = in0;
    end

    reg [7:0] out2119;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2119 = in0;
    end

    reg [7:0] out2120;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2120 = in0;
    end

    reg [7:0] out2121;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2121 = in0;
    end

    reg [7:0] out2122;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2122 = in0;
    end

    reg [7:0] out2123;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2123 = in0;
    end

    reg [7:0] out2124;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2124 = in0;
    end

    reg [7:0] out2125;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2125 = in0;
    end

    reg [7:0] out2126;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2126 = in0;
    end

    reg [7:0] out2127;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2127 = in0;
    end

    reg [7:0] out2128;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2128 = in0;
    end

    reg [7:0] out2129;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2129 = in0;
    end

    reg [7:0] out2130;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2130 = in0;
    end

    reg [7:0] out2131;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2131 = in0;
    end

    reg [7:0] out2132;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2132 = in0;
    end

    reg [7:0] out2133;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2133 = in0;
    end

    reg [7:0] out2134;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2134 = in0;
    end

    reg [7:0] out2135;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2135 = in0;
    end

    reg [7:0] out2136;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2136 = in0;
    end

    reg [7:0] out2137;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2137 = in0;
    end

    reg [7:0] out2138;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2138 = in0;
    end

    reg [7:0] out2139;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2139 = in0;
    end

    reg [7:0] out2140;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2140 = in0;
    end

    reg [7:0] out2141;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2141 = in0;
    end

    reg [7:0] out2142;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2142 = in0;
    end

    reg [7:0] out2143;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2143 = in0;
    end

    reg [7:0] out2144;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2144 = in0;
    end

    reg [7:0] out2145;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2145 = in0;
    end

    reg [7:0] out2146;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2146 = in0;
    end

    reg [7:0] out2147;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2147 = in0;
    end

    reg [7:0] out2148;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2148 = in0;
    end

    reg [7:0] out2149;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2149 = in0;
    end

    reg [7:0] out2150;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2150 = in0;
    end

    reg [7:0] out2151;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2151 = in0;
    end

    reg [7:0] out2152;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2152 = in0;
    end

    reg [7:0] out2153;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2153 = in0;
    end

    reg [7:0] out2154;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2154 = in0;
    end

    reg [7:0] out2155;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2155 = in0;
    end

    reg [7:0] out2156;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2156 = in0;
    end

    reg [7:0] out2157;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2157 = in0;
    end

    reg [7:0] out2158;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2158 = in0;
    end

    reg [7:0] out2159;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2159 = in0;
    end

    reg [7:0] out2160;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2160 = in0;
    end

    reg [7:0] out2161;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2161 = in0;
    end

    reg [7:0] out2162;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2162 = in0;
    end

    reg [7:0] out2163;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2163 = in0;
    end

    reg [7:0] out2164;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2164 = in0;
    end

    reg [7:0] out2165;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2165 = in0;
    end

    reg [7:0] out2166;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2166 = in0;
    end

    reg [7:0] out2167;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2167 = in0;
    end

    reg [7:0] out2168;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2168 = in0;
    end

    reg [7:0] out2169;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2169 = in0;
    end

    reg [7:0] out2170;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2170 = in0;
    end

    reg [7:0] out2171;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2171 = in0;
    end

    reg [7:0] out2172;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2172 = in0;
    end

    reg [7:0] out2173;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2173 = in0;
    end

    reg [7:0] out2174;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2174 = in0;
    end

    reg [7:0] out2175;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2175 = in0;
    end

    reg [7:0] out2176;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2176 = in0;
    end

    reg [7:0] out2177;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2177 = in0;
    end

    reg [7:0] out2178;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2178 = in0;
    end

    reg [7:0] out2179;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2179 = in0;
    end

    reg [7:0] out2180;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2180 = in0;
    end

    reg [7:0] out2181;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2181 = in0;
    end

    reg [7:0] out2182;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2182 = in0;
    end

    reg [7:0] out2183;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2183 = in0;
    end

    reg [7:0] out2184;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2184 = in0;
    end

    reg [7:0] out2185;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2185 = in0;
    end

    reg [7:0] out2186;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2186 = in0;
    end

    reg [7:0] out2187;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2187 = in0;
    end

    reg [7:0] out2188;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2188 = in0;
    end

    reg [7:0] out2189;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2189 = in0;
    end

    reg [7:0] out2190;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2190 = in0;
    end

    reg [7:0] out2191;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2191 = in0;
    end

    reg [7:0] out2192;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2192 = in0;
    end

    reg [7:0] out2193;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2193 = in0;
    end

    reg [7:0] out2194;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2194 = in0;
    end

    reg [7:0] out2195;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2195 = in0;
    end

    reg [7:0] out2196;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2196 = in0;
    end

    reg [7:0] out2197;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2197 = in0;
    end

    reg [7:0] out2198;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2198 = in0;
    end

    reg [7:0] out2199;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2199 = in0;
    end

    reg [7:0] out2200;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2200 = in0;
    end

    reg [7:0] out2201;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2201 = in0;
    end

    reg [7:0] out2202;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2202 = in0;
    end

    reg [7:0] out2203;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2203 = in0;
    end

    reg [7:0] out2204;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2204 = in0;
    end

    reg [7:0] out2205;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2205 = in0;
    end

    reg [7:0] out2206;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2206 = in0;
    end

    reg [7:0] out2207;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2207 = in0;
    end

    reg [7:0] out2208;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2208 = in0;
    end

    reg [7:0] out2209;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2209 = in0;
    end

    reg [7:0] out2210;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2210 = in0;
    end

    reg [7:0] out2211;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2211 = in0;
    end

    reg [7:0] out2212;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2212 = in0;
    end

    reg [7:0] out2213;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2213 = in0;
    end

    reg [7:0] out2214;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2214 = in0;
    end

    reg [7:0] out2215;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2215 = in0;
    end

    reg [7:0] out2216;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2216 = in0;
    end

    reg [7:0] out2217;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2217 = in0;
    end

    reg [7:0] out2218;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2218 = in0;
    end

    reg [7:0] out2219;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2219 = in0;
    end

    reg [7:0] out2220;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2220 = in0;
    end

    reg [7:0] out2221;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2221 = in0;
    end

    reg [7:0] out2222;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2222 = in0;
    end

    reg [7:0] out2223;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2223 = in0;
    end

    reg [7:0] out2224;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2224 = in0;
    end

    reg [7:0] out2225;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2225 = in0;
    end

    reg [7:0] out2226;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2226 = in0;
    end

    reg [7:0] out2227;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2227 = in0;
    end

    reg [7:0] out2228;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2228 = in0;
    end

    reg [7:0] out2229;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2229 = in0;
    end

    reg [7:0] out2230;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2230 = in0;
    end

    reg [7:0] out2231;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2231 = in0;
    end

    reg [7:0] out2232;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2232 = in0;
    end

    reg [7:0] out2233;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2233 = in0;
    end

    reg [7:0] out2234;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2234 = in0;
    end

    reg [7:0] out2235;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2235 = in0;
    end

    reg [7:0] out2236;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2236 = in0;
    end

    reg [7:0] out2237;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2237 = in0;
    end

    reg [7:0] out2238;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2238 = in0;
    end

    reg [7:0] out2239;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2239 = in0;
    end

    reg [7:0] out2240;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2240 = in0;
    end

    reg [7:0] out2241;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2241 = in0;
    end

    reg [7:0] out2242;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2242 = in0;
    end

    reg [7:0] out2243;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2243 = in0;
    end

    reg [7:0] out2244;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2244 = in0;
    end

    reg [7:0] out2245;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2245 = in0;
    end

    reg [7:0] out2246;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2246 = in0;
    end

    reg [7:0] out2247;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2247 = in0;
    end

    reg [7:0] out2248;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2248 = in0;
    end

    reg [7:0] out2249;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2249 = in0;
    end

    reg [7:0] out2250;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2250 = in0;
    end

    reg [7:0] out2251;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2251 = in0;
    end

    reg [7:0] out2252;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2252 = in0;
    end

    reg [7:0] out2253;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2253 = in0;
    end

    reg [7:0] out2254;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2254 = in0;
    end

    reg [7:0] out2255;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2255 = in0;
    end

    reg [7:0] out2256;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2256 = in0;
    end

    reg [7:0] out2257;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2257 = in0;
    end

    reg [7:0] out2258;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2258 = in0;
    end

    reg [7:0] out2259;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2259 = in0;
    end

    reg [7:0] out2260;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2260 = in0;
    end

    reg [7:0] out2261;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2261 = in0;
    end

    reg [7:0] out2262;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2262 = in0;
    end

    reg [7:0] out2263;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2263 = in0;
    end

    reg [7:0] out2264;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2264 = in0;
    end

    reg [7:0] out2265;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2265 = in0;
    end

    reg [7:0] out2266;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2266 = in0;
    end

    reg [7:0] out2267;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2267 = in0;
    end

    reg [7:0] out2268;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2268 = in0;
    end

    reg [7:0] out2269;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2269 = in0;
    end

    reg [7:0] out2270;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2270 = in0;
    end

    reg [7:0] out2271;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2271 = in0;
    end

    reg [7:0] out2272;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2272 = in0;
    end

    reg [7:0] out2273;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2273 = in0;
    end

    reg [7:0] out2274;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2274 = in0;
    end

    reg [7:0] out2275;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2275 = in0;
    end

    reg [7:0] out2276;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2276 = in0;
    end

    reg [7:0] out2277;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2277 = in0;
    end

    reg [7:0] out2278;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2278 = in0;
    end

    reg [7:0] out2279;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2279 = in0;
    end

    reg [7:0] out2280;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2280 = in0;
    end

    reg [7:0] out2281;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2281 = in0;
    end

    reg [7:0] out2282;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2282 = in0;
    end

    reg [7:0] out2283;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2283 = in0;
    end

    reg [7:0] out2284;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2284 = in0;
    end

    reg [7:0] out2285;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2285 = in0;
    end

    reg [7:0] out2286;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2286 = in0;
    end

    reg [7:0] out2287;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2287 = in0;
    end

    reg [7:0] out2288;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2288 = in0;
    end

    reg [7:0] out2289;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2289 = in0;
    end

    reg [7:0] out2290;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2290 = in0;
    end

    reg [7:0] out2291;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2291 = in0;
    end

    reg [7:0] out2292;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2292 = in0;
    end

    reg [7:0] out2293;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2293 = in0;
    end

    reg [7:0] out2294;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2294 = in0;
    end

    reg [7:0] out2295;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2295 = in0;
    end

    reg [7:0] out2296;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2296 = in0;
    end

    reg [7:0] out2297;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2297 = in0;
    end

    reg [7:0] out2298;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2298 = in0;
    end

    reg [7:0] out2299;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2299 = in0;
    end

    reg [7:0] out2300;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2300 = in0;
    end

    reg [7:0] out2301;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2301 = in0;
    end

    reg [7:0] out2302;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2302 = in0;
    end

    reg [7:0] out2303;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2303 = in0;
    end

    reg [7:0] out2304;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2304 = in0;
    end

    reg [7:0] out2305;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2305 = in0;
    end

    reg [7:0] out2306;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2306 = in0;
    end

    reg [7:0] out2307;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2307 = in0;
    end

    reg [7:0] out2308;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2308 = in0;
    end

    reg [7:0] out2309;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2309 = in0;
    end

    reg [7:0] out2310;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2310 = in0;
    end

    reg [7:0] out2311;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2311 = in0;
    end

    reg [7:0] out2312;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2312 = in0;
    end

    reg [7:0] out2313;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2313 = in0;
    end

    reg [7:0] out2314;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2314 = in0;
    end

    reg [7:0] out2315;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2315 = in0;
    end

    reg [7:0] out2316;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2316 = in0;
    end

    reg [7:0] out2317;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2317 = in0;
    end

    reg [7:0] out2318;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2318 = in0;
    end

    reg [7:0] out2319;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2319 = in0;
    end

    reg [7:0] out2320;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2320 = in0;
    end

    reg [7:0] out2321;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2321 = in0;
    end

    reg [7:0] out2322;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2322 = in0;
    end

    reg [7:0] out2323;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2323 = in0;
    end

    reg [7:0] out2324;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2324 = in0;
    end

    reg [7:0] out2325;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2325 = in0;
    end

    reg [7:0] out2326;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2326 = in0;
    end

    reg [7:0] out2327;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2327 = in0;
    end

    reg [7:0] out2328;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2328 = in0;
    end

    reg [7:0] out2329;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2329 = in0;
    end

    reg [7:0] out2330;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2330 = in0;
    end

    reg [7:0] out2331;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2331 = in0;
    end

    reg [7:0] out2332;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2332 = in0;
    end

    reg [7:0] out2333;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2333 = in0;
    end

    reg [7:0] out2334;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2334 = in0;
    end

    reg [7:0] out2335;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2335 = in0;
    end

    reg [7:0] out2336;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2336 = in0;
    end

    reg [7:0] out2337;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2337 = in0;
    end

    reg [7:0] out2338;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2338 = in0;
    end

    reg [7:0] out2339;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2339 = in0;
    end

    reg [7:0] out2340;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2340 = in0;
    end

    reg [7:0] out2341;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2341 = in0;
    end

    reg [7:0] out2342;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2342 = in0;
    end

    reg [7:0] out2343;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2343 = in0;
    end

    reg [7:0] out2344;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2344 = in0;
    end

    reg [7:0] out2345;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2345 = in0;
    end

    reg [7:0] out2346;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2346 = in0;
    end

    reg [7:0] out2347;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2347 = in0;
    end

    reg [7:0] out2348;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2348 = in0;
    end

    reg [7:0] out2349;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2349 = in0;
    end

    reg [7:0] out2350;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2350 = in0;
    end

    reg [7:0] out2351;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2351 = in0;
    end

    reg [7:0] out2352;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2352 = in0;
    end

    reg [7:0] out2353;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2353 = in0;
    end

    reg [7:0] out2354;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2354 = in0;
    end

    reg [7:0] out2355;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2355 = in0;
    end

    reg [7:0] out2356;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2356 = in0;
    end

    reg [7:0] out2357;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2357 = in0;
    end

    reg [7:0] out2358;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2358 = in0;
    end

    reg [7:0] out2359;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2359 = in0;
    end

    reg [7:0] out2360;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2360 = in0;
    end

    reg [7:0] out2361;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2361 = in0;
    end

    reg [7:0] out2362;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2362 = in0;
    end

    reg [7:0] out2363;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2363 = in0;
    end

    reg [7:0] out2364;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2364 = in0;
    end

    reg [7:0] out2365;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2365 = in0;
    end

    reg [7:0] out2366;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2366 = in0;
    end

    reg [7:0] out2367;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2367 = in0;
    end

    reg [7:0] out2368;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2368 = in0;
    end

    reg [7:0] out2369;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2369 = in0;
    end

    reg [7:0] out2370;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2370 = in0;
    end

    reg [7:0] out2371;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2371 = in0;
    end

    reg [7:0] out2372;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2372 = in0;
    end

    reg [7:0] out2373;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2373 = in0;
    end

    reg [7:0] out2374;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2374 = in0;
    end

    reg [7:0] out2375;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2375 = in0;
    end

    reg [7:0] out2376;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2376 = in0;
    end

    reg [7:0] out2377;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2377 = in0;
    end

    reg [7:0] out2378;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2378 = in0;
    end

    reg [7:0] out2379;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2379 = in0;
    end

    reg [7:0] out2380;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2380 = in0;
    end

    reg [7:0] out2381;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2381 = in0;
    end

    reg [7:0] out2382;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2382 = in0;
    end

    reg [7:0] out2383;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2383 = in0;
    end

    reg [7:0] out2384;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2384 = in0;
    end

    reg [7:0] out2385;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2385 = in0;
    end

    reg [7:0] out2386;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2386 = in0;
    end

    reg [7:0] out2387;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2387 = in0;
    end

    reg [7:0] out2388;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2388 = in0;
    end

    reg [7:0] out2389;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2389 = in0;
    end

    reg [7:0] out2390;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2390 = in0;
    end

    reg [7:0] out2391;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2391 = in0;
    end

    reg [7:0] out2392;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2392 = in0;
    end

    reg [7:0] out2393;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2393 = in0;
    end

    reg [7:0] out2394;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2394 = in0;
    end

    reg [7:0] out2395;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2395 = in0;
    end

    reg [7:0] out2396;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2396 = in0;
    end

    reg [7:0] out2397;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2397 = in0;
    end

    reg [7:0] out2398;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2398 = in0;
    end

    reg [7:0] out2399;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2399 = in0;
    end

    reg [7:0] out2400;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2400 = in0;
    end

    reg [7:0] out2401;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2401 = in0;
    end

    reg [7:0] out2402;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2402 = in0;
    end

    reg [7:0] out2403;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2403 = in0;
    end

    reg [7:0] out2404;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2404 = in0;
    end

    reg [7:0] out2405;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2405 = in0;
    end

    reg [7:0] out2406;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2406 = in0;
    end

    reg [7:0] out2407;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2407 = in0;
    end

    reg [7:0] out2408;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2408 = in0;
    end

    reg [7:0] out2409;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2409 = in0;
    end

    reg [7:0] out2410;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2410 = in0;
    end

    reg [7:0] out2411;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2411 = in0;
    end

    reg [7:0] out2412;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2412 = in0;
    end

    reg [7:0] out2413;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2413 = in0;
    end

    reg [7:0] out2414;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2414 = in0;
    end

    reg [7:0] out2415;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2415 = in0;
    end

    reg [7:0] out2416;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2416 = in0;
    end

    reg [7:0] out2417;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2417 = in0;
    end

    reg [7:0] out2418;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2418 = in0;
    end

    reg [7:0] out2419;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2419 = in0;
    end

    reg [7:0] out2420;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2420 = in0;
    end

    reg [7:0] out2421;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2421 = in0;
    end

    reg [7:0] out2422;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2422 = in0;
    end

    reg [7:0] out2423;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2423 = in0;
    end

    reg [7:0] out2424;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2424 = in0;
    end

    reg [7:0] out2425;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2425 = in0;
    end

    reg [7:0] out2426;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2426 = in0;
    end

    reg [7:0] out2427;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2427 = in0;
    end

    reg [7:0] out2428;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2428 = in0;
    end

    reg [7:0] out2429;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2429 = in0;
    end

    reg [7:0] out2430;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2430 = in0;
    end

    reg [7:0] out2431;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2431 = in0;
    end

    reg [7:0] out2432;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2432 = in0;
    end

    reg [7:0] out2433;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2433 = in0;
    end

    reg [7:0] out2434;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2434 = in0;
    end

    reg [7:0] out2435;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2435 = in0;
    end

    reg [7:0] out2436;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2436 = in0;
    end

    reg [7:0] out2437;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2437 = in0;
    end

    reg [7:0] out2438;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2438 = in0;
    end

    reg [7:0] out2439;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2439 = in0;
    end

    reg [7:0] out2440;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2440 = in0;
    end

    reg [7:0] out2441;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2441 = in0;
    end

    reg [7:0] out2442;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2442 = in0;
    end

    reg [7:0] out2443;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2443 = in0;
    end

    reg [7:0] out2444;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2444 = in0;
    end

    reg [7:0] out2445;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2445 = in0;
    end

    reg [7:0] out2446;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2446 = in0;
    end

    reg [7:0] out2447;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2447 = in0;
    end

    reg [7:0] out2448;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2448 = in0;
    end

    reg [7:0] out2449;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2449 = in0;
    end

    reg [7:0] out2450;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2450 = in0;
    end

    reg [7:0] out2451;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2451 = in0;
    end

    reg [7:0] out2452;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2452 = in0;
    end

    reg [7:0] out2453;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2453 = in0;
    end

    reg [7:0] out2454;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2454 = in0;
    end

    reg [7:0] out2455;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2455 = in0;
    end

    reg [7:0] out2456;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2456 = in0;
    end

    reg [7:0] out2457;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2457 = in0;
    end

    reg [7:0] out2458;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2458 = in0;
    end

    reg [7:0] out2459;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2459 = in0;
    end

    reg [7:0] out2460;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2460 = in0;
    end

    reg [7:0] out2461;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2461 = in0;
    end

    reg [7:0] out2462;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2462 = in0;
    end

    reg [7:0] out2463;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2463 = in0;
    end

    reg [7:0] out2464;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2464 = in0;
    end

    reg [7:0] out2465;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2465 = in0;
    end

    reg [7:0] out2466;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2466 = in0;
    end

    reg [7:0] out2467;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2467 = in0;
    end

    reg [7:0] out2468;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2468 = in0;
    end

    reg [7:0] out2469;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2469 = in0;
    end

    reg [7:0] out2470;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2470 = in0;
    end

    reg [7:0] out2471;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2471 = in0;
    end

    reg [7:0] out2472;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2472 = in0;
    end

    reg [7:0] out2473;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2473 = in0;
    end

    reg [7:0] out2474;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2474 = in0;
    end

    reg [7:0] out2475;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2475 = in0;
    end

    reg [7:0] out2476;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2476 = in0;
    end

    reg [7:0] out2477;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2477 = in0;
    end

    reg [7:0] out2478;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2478 = in0;
    end

    reg [7:0] out2479;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2479 = in0;
    end

    reg [7:0] out2480;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2480 = in0;
    end

    reg [7:0] out2481;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2481 = in0;
    end

    reg [7:0] out2482;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2482 = in0;
    end

    reg [7:0] out2483;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2483 = in0;
    end

    reg [7:0] out2484;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2484 = in0;
    end

    reg [7:0] out2485;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2485 = in0;
    end

    reg [7:0] out2486;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2486 = in0;
    end

    reg [7:0] out2487;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2487 = in0;
    end

    reg [7:0] out2488;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2488 = in0;
    end

    reg [7:0] out2489;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2489 = in0;
    end

    reg [7:0] out2490;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2490 = in0;
    end

    reg [7:0] out2491;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2491 = in0;
    end

    reg [7:0] out2492;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2492 = in0;
    end

    reg [7:0] out2493;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2493 = in0;
    end

    reg [7:0] out2494;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2494 = in0;
    end

    reg [7:0] out2495;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2495 = in0;
    end

    reg [7:0] out2496;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2496 = in0;
    end

    reg [7:0] out2497;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2497 = in0;
    end

    reg [7:0] out2498;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2498 = in0;
    end

    reg [7:0] out2499;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2499 = in0;
    end

    reg [7:0] out2500;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2500 = in0;
    end

    reg [7:0] out2501;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2501 = in0;
    end

    reg [7:0] out2502;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2502 = in0;
    end

    reg [7:0] out2503;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2503 = in0;
    end

    reg [7:0] out2504;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2504 = in0;
    end

    reg [7:0] out2505;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2505 = in0;
    end

    reg [7:0] out2506;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2506 = in0;
    end

    reg [7:0] out2507;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2507 = in0;
    end

    reg [7:0] out2508;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2508 = in0;
    end

    reg [7:0] out2509;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2509 = in0;
    end

    reg [7:0] out2510;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2510 = in0;
    end

    reg [7:0] out2511;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2511 = in0;
    end

    reg [7:0] out2512;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2512 = in0;
    end

    reg [7:0] out2513;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2513 = in0;
    end

    reg [7:0] out2514;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2514 = in0;
    end

    reg [7:0] out2515;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2515 = in0;
    end

    reg [7:0] out2516;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2516 = in0;
    end

    reg [7:0] out2517;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2517 = in0;
    end

    reg [7:0] out2518;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2518 = in0;
    end

    reg [7:0] out2519;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2519 = in0;
    end

    reg [7:0] out2520;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2520 = in0;
    end

    reg [7:0] out2521;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2521 = in0;
    end

    reg [7:0] out2522;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2522 = in0;
    end

    reg [7:0] out2523;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2523 = in0;
    end

    reg [7:0] out2524;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2524 = in0;
    end

    reg [7:0] out2525;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2525 = in0;
    end

    reg [7:0] out2526;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2526 = in0;
    end

    reg [7:0] out2527;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2527 = in0;
    end

    reg [7:0] out2528;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2528 = in0;
    end

    reg [7:0] out2529;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2529 = in0;
    end

    reg [7:0] out2530;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2530 = in0;
    end

    reg [7:0] out2531;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2531 = in0;
    end

    reg [7:0] out2532;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2532 = in0;
    end

    reg [7:0] out2533;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2533 = in0;
    end

    reg [7:0] out2534;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2534 = in0;
    end

    reg [7:0] out2535;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2535 = in0;
    end

    reg [7:0] out2536;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2536 = in0;
    end

    reg [7:0] out2537;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2537 = in0;
    end

    reg [7:0] out2538;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2538 = in0;
    end

    reg [7:0] out2539;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2539 = in0;
    end

    reg [7:0] out2540;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2540 = in0;
    end

    reg [7:0] out2541;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2541 = in0;
    end

    reg [7:0] out2542;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2542 = in0;
    end

    reg [7:0] out2543;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2543 = in0;
    end

    reg [7:0] out2544;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2544 = in0;
    end

    reg [7:0] out2545;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2545 = in0;
    end

    reg [7:0] out2546;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2546 = in0;
    end

    reg [7:0] out2547;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2547 = in0;
    end

    reg [7:0] out2548;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2548 = in0;
    end

    reg [7:0] out2549;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2549 = in0;
    end

    reg [7:0] out2550;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2550 = in0;
    end

    reg [7:0] out2551;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2551 = in0;
    end

    reg [7:0] out2552;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2552 = in0;
    end

    reg [7:0] out2553;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2553 = in0;
    end

    reg [7:0] out2554;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2554 = in0;
    end

    reg [7:0] out2555;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2555 = in0;
    end

    reg [7:0] out2556;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2556 = in0;
    end

    reg [7:0] out2557;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2557 = in0;
    end

    reg [7:0] out2558;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2558 = in0;
    end

    reg [7:0] out2559;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2559 = in0;
    end

    reg [7:0] out2560;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2560 = in0;
    end

    reg [7:0] out2561;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2561 = in0;
    end

    reg [7:0] out2562;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2562 = in0;
    end

    reg [7:0] out2563;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2563 = in0;
    end

    reg [7:0] out2564;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2564 = in0;
    end

    reg [7:0] out2565;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2565 = in0;
    end

    reg [7:0] out2566;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2566 = in0;
    end

    reg [7:0] out2567;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2567 = in0;
    end

    reg [7:0] out2568;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2568 = in0;
    end

    reg [7:0] out2569;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2569 = in0;
    end

    reg [7:0] out2570;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2570 = in0;
    end

    reg [7:0] out2571;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2571 = in0;
    end

    reg [7:0] out2572;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2572 = in0;
    end

    reg [7:0] out2573;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2573 = in0;
    end

    reg [7:0] out2574;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2574 = in0;
    end

    reg [7:0] out2575;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2575 = in0;
    end

    reg [7:0] out2576;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2576 = in0;
    end

    reg [7:0] out2577;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2577 = in0;
    end

    reg [7:0] out2578;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2578 = in0;
    end

    reg [7:0] out2579;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2579 = in0;
    end

    reg [7:0] out2580;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2580 = in0;
    end

    reg [7:0] out2581;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2581 = in0;
    end

    reg [7:0] out2582;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2582 = in0;
    end

    reg [7:0] out2583;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2583 = in0;
    end

    reg [7:0] out2584;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2584 = in0;
    end

    reg [7:0] out2585;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2585 = in0;
    end

    reg [7:0] out2586;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2586 = in0;
    end

    reg [7:0] out2587;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2587 = in0;
    end

    reg [7:0] out2588;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2588 = in0;
    end

    reg [7:0] out2589;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2589 = in0;
    end

    reg [7:0] out2590;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2590 = in0;
    end

    reg [7:0] out2591;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2591 = in0;
    end

    reg [7:0] out2592;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2592 = in0;
    end

    reg [7:0] out2593;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2593 = in0;
    end

    reg [7:0] out2594;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2594 = in0;
    end

    reg [7:0] out2595;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2595 = in0;
    end

    reg [7:0] out2596;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2596 = in0;
    end

    reg [7:0] out2597;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2597 = in0;
    end

    reg [7:0] out2598;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2598 = in0;
    end

    reg [7:0] out2599;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2599 = in0;
    end

    reg [7:0] out2600;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2600 = in0;
    end

    reg [7:0] out2601;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2601 = in0;
    end

    reg [7:0] out2602;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2602 = in0;
    end

    reg [7:0] out2603;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2603 = in0;
    end

    reg [7:0] out2604;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2604 = in0;
    end

    reg [7:0] out2605;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2605 = in0;
    end

    reg [7:0] out2606;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2606 = in0;
    end

    reg [7:0] out2607;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2607 = in0;
    end

    reg [7:0] out2608;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2608 = in0;
    end

    reg [7:0] out2609;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2609 = in0;
    end

    reg [7:0] out2610;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2610 = in0;
    end

    reg [7:0] out2611;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2611 = in0;
    end

    reg [7:0] out2612;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2612 = in0;
    end

    reg [7:0] out2613;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2613 = in0;
    end

    reg [7:0] out2614;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2614 = in0;
    end

    reg [7:0] out2615;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2615 = in0;
    end

    reg [7:0] out2616;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2616 = in0;
    end

    reg [7:0] out2617;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2617 = in0;
    end

    reg [7:0] out2618;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2618 = in0;
    end

    reg [7:0] out2619;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2619 = in0;
    end

    reg [7:0] out2620;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2620 = in0;
    end

    reg [7:0] out2621;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2621 = in0;
    end

    reg [7:0] out2622;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2622 = in0;
    end

    reg [7:0] out2623;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2623 = in0;
    end

    reg [7:0] out2624;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2624 = in0;
    end

    reg [7:0] out2625;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2625 = in0;
    end

    reg [7:0] out2626;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2626 = in0;
    end

    reg [7:0] out2627;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2627 = in0;
    end

    reg [7:0] out2628;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2628 = in0;
    end

    reg [7:0] out2629;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2629 = in0;
    end

    reg [7:0] out2630;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2630 = in0;
    end

    reg [7:0] out2631;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2631 = in0;
    end

    reg [7:0] out2632;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2632 = in0;
    end

    reg [7:0] out2633;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2633 = in0;
    end

    reg [7:0] out2634;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2634 = in0;
    end

    reg [7:0] out2635;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2635 = in0;
    end

    reg [7:0] out2636;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2636 = in0;
    end

    reg [7:0] out2637;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2637 = in0;
    end

    reg [7:0] out2638;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2638 = in0;
    end

    reg [7:0] out2639;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2639 = in0;
    end

    reg [7:0] out2640;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2640 = in0;
    end

    reg [7:0] out2641;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2641 = in0;
    end

    reg [7:0] out2642;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2642 = in0;
    end

    reg [7:0] out2643;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2643 = in0;
    end

    reg [7:0] out2644;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2644 = in0;
    end

    reg [7:0] out2645;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2645 = in0;
    end

    reg [7:0] out2646;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2646 = in0;
    end

    reg [7:0] out2647;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2647 = in0;
    end

    reg [7:0] out2648;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2648 = in0;
    end

    reg [7:0] out2649;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2649 = in0;
    end

    reg [7:0] out2650;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2650 = in0;
    end

    reg [7:0] out2651;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2651 = in0;
    end

    reg [7:0] out2652;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2652 = in0;
    end

    reg [7:0] out2653;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2653 = in0;
    end

    reg [7:0] out2654;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2654 = in0;
    end

    reg [7:0] out2655;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2655 = in0;
    end

    reg [7:0] out2656;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2656 = in0;
    end

    reg [7:0] out2657;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2657 = in0;
    end

    reg [7:0] out2658;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2658 = in0;
    end

    reg [7:0] out2659;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2659 = in0;
    end

    reg [7:0] out2660;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2660 = in0;
    end

    reg [7:0] out2661;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2661 = in0;
    end

    reg [7:0] out2662;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2662 = in0;
    end

    reg [7:0] out2663;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2663 = in0;
    end

    reg [7:0] out2664;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2664 = in0;
    end

    reg [7:0] out2665;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2665 = in0;
    end

    reg [7:0] out2666;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2666 = in0;
    end

    reg [7:0] out2667;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2667 = in0;
    end

    reg [7:0] out2668;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2668 = in0;
    end

    reg [7:0] out2669;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2669 = in0;
    end

    reg [7:0] out2670;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2670 = in0;
    end

    reg [7:0] out2671;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2671 = in0;
    end

    reg [7:0] out2672;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2672 = in0;
    end

    reg [7:0] out2673;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2673 = in0;
    end

    reg [7:0] out2674;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2674 = in0;
    end

    reg [7:0] out2675;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2675 = in0;
    end

    reg [7:0] out2676;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2676 = in0;
    end

    reg [7:0] out2677;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2677 = in0;
    end

    reg [7:0] out2678;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2678 = in0;
    end

    reg [7:0] out2679;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2679 = in0;
    end

    reg [7:0] out2680;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2680 = in0;
    end

    reg [7:0] out2681;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2681 = in0;
    end

    reg [7:0] out2682;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2682 = in0;
    end

    reg [7:0] out2683;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2683 = in0;
    end

    reg [7:0] out2684;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2684 = in0;
    end

    reg [7:0] out2685;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2685 = in0;
    end

    reg [7:0] out2686;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2686 = in0;
    end

    reg [7:0] out2687;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2687 = in0;
    end

    reg [7:0] out2688;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2688 = in0;
    end

    reg [7:0] out2689;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2689 = in0;
    end

    reg [7:0] out2690;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2690 = in0;
    end

    reg [7:0] out2691;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2691 = in0;
    end

    reg [7:0] out2692;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2692 = in0;
    end

    reg [7:0] out2693;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2693 = in0;
    end

    reg [7:0] out2694;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2694 = in0;
    end

    reg [7:0] out2695;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2695 = in0;
    end

    reg [7:0] out2696;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2696 = in0;
    end

    reg [7:0] out2697;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2697 = in0;
    end

    reg [7:0] out2698;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2698 = in0;
    end

    reg [7:0] out2699;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2699 = in0;
    end

    reg [7:0] out2700;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2700 = in0;
    end

    reg [7:0] out2701;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2701 = in0;
    end

    reg [7:0] out2702;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2702 = in0;
    end

    reg [7:0] out2703;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2703 = in0;
    end

    reg [7:0] out2704;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2704 = in0;
    end

    reg [7:0] out2705;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2705 = in0;
    end

    reg [7:0] out2706;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2706 = in0;
    end

    reg [7:0] out2707;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2707 = in0;
    end

    reg [7:0] out2708;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2708 = in0;
    end

    reg [7:0] out2709;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2709 = in0;
    end

    reg [7:0] out2710;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2710 = in0;
    end

    reg [7:0] out2711;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2711 = in0;
    end

    reg [7:0] out2712;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2712 = in0;
    end

    reg [7:0] out2713;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2713 = in0;
    end

    reg [7:0] out2714;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2714 = in0;
    end

    reg [7:0] out2715;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2715 = in0;
    end

    reg [7:0] out2716;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2716 = in0;
    end

    reg [7:0] out2717;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2717 = in0;
    end

    reg [7:0] out2718;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2718 = in0;
    end

    reg [7:0] out2719;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2719 = in0;
    end

    reg [7:0] out2720;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2720 = in0;
    end

    reg [7:0] out2721;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2721 = in0;
    end

    reg [7:0] out2722;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2722 = in0;
    end

    reg [7:0] out2723;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2723 = in0;
    end

    reg [7:0] out2724;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2724 = in0;
    end

    reg [7:0] out2725;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2725 = in0;
    end

    reg [7:0] out2726;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2726 = in0;
    end

    reg [7:0] out2727;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2727 = in0;
    end

    reg [7:0] out2728;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2728 = in0;
    end

    reg [7:0] out2729;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2729 = in0;
    end

    reg [7:0] out2730;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2730 = in0;
    end

    reg [7:0] out2731;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2731 = in0;
    end

    reg [7:0] out2732;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2732 = in0;
    end

    reg [7:0] out2733;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2733 = in0;
    end

    reg [7:0] out2734;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2734 = in0;
    end

    reg [7:0] out2735;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2735 = in0;
    end

    reg [7:0] out2736;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2736 = in0;
    end

    reg [7:0] out2737;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2737 = in0;
    end

    reg [7:0] out2738;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2738 = in0;
    end

    reg [7:0] out2739;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2739 = in0;
    end

    reg [7:0] out2740;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2740 = in0;
    end

    reg [7:0] out2741;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2741 = in0;
    end

    reg [7:0] out2742;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2742 = in0;
    end

    reg [7:0] out2743;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2743 = in0;
    end

    reg [7:0] out2744;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2744 = in0;
    end

    reg [7:0] out2745;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2745 = in0;
    end

    reg [7:0] out2746;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2746 = in0;
    end

    reg [7:0] out2747;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2747 = in0;
    end

    reg [7:0] out2748;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2748 = in0;
    end

    reg [7:0] out2749;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2749 = in0;
    end

    reg [7:0] out2750;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2750 = in0;
    end

    reg [7:0] out2751;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2751 = in0;
    end

    reg [7:0] out2752;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2752 = in0;
    end

    reg [7:0] out2753;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2753 = in0;
    end

    reg [7:0] out2754;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2754 = in0;
    end

    reg [7:0] out2755;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2755 = in0;
    end

    reg [7:0] out2756;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2756 = in0;
    end

    reg [7:0] out2757;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2757 = in0;
    end

    reg [7:0] out2758;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2758 = in0;
    end

    reg [7:0] out2759;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2759 = in0;
    end

    reg [7:0] out2760;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2760 = in0;
    end

    reg [7:0] out2761;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2761 = in0;
    end

    reg [7:0] out2762;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2762 = in0;
    end

    reg [7:0] out2763;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2763 = in0;
    end

    reg [7:0] out2764;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2764 = in0;
    end

    reg [7:0] out2765;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2765 = in0;
    end

    reg [7:0] out2766;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2766 = in0;
    end

    reg [7:0] out2767;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2767 = in0;
    end

    reg [7:0] out2768;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2768 = in0;
    end

    reg [7:0] out2769;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2769 = in0;
    end

    reg [7:0] out2770;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2770 = in0;
    end

    reg [7:0] out2771;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2771 = in0;
    end

    reg [7:0] out2772;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2772 = in0;
    end

    reg [7:0] out2773;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2773 = in0;
    end

    reg [7:0] out2774;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2774 = in0;
    end

    reg [7:0] out2775;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2775 = in0;
    end

    reg [7:0] out2776;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2776 = in0;
    end

    reg [7:0] out2777;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2777 = in0;
    end

    reg [7:0] out2778;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2778 = in0;
    end

    reg [7:0] out2779;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2779 = in0;
    end

    reg [7:0] out2780;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2780 = in0;
    end

    reg [7:0] out2781;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2781 = in0;
    end

    reg [7:0] out2782;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2782 = in0;
    end

    reg [7:0] out2783;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2783 = in0;
    end

    reg [7:0] out2784;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2784 = in0;
    end

    reg [7:0] out2785;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2785 = in0;
    end

    reg [7:0] out2786;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2786 = in0;
    end

    reg [7:0] out2787;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2787 = in0;
    end

    reg [7:0] out2788;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2788 = in0;
    end

    reg [7:0] out2789;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2789 = in0;
    end

    reg [7:0] out2790;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2790 = in0;
    end

    reg [7:0] out2791;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2791 = in0;
    end

    reg [7:0] out2792;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2792 = in0;
    end

    reg [7:0] out2793;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2793 = in0;
    end

    reg [7:0] out2794;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2794 = in0;
    end

    reg [7:0] out2795;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2795 = in0;
    end

    reg [7:0] out2796;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2796 = in0;
    end

    reg [7:0] out2797;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2797 = in0;
    end

    reg [7:0] out2798;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2798 = in0;
    end

    reg [7:0] out2799;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2799 = in0;
    end

    reg [7:0] out2800;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2800 = in0;
    end

    reg [7:0] out2801;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2801 = in0;
    end

    reg [7:0] out2802;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2802 = in0;
    end

    reg [7:0] out2803;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2803 = in0;
    end

    reg [7:0] out2804;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2804 = in0;
    end

    reg [7:0] out2805;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2805 = in0;
    end

    reg [7:0] out2806;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2806 = in0;
    end

    reg [7:0] out2807;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2807 = in0;
    end

    reg [7:0] out2808;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2808 = in0;
    end

    reg [7:0] out2809;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2809 = in0;
    end

    reg [7:0] out2810;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2810 = in0;
    end

    reg [7:0] out2811;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2811 = in0;
    end

    reg [7:0] out2812;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2812 = in0;
    end

    reg [7:0] out2813;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2813 = in0;
    end

    reg [7:0] out2814;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2814 = in0;
    end

    reg [7:0] out2815;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2815 = in0;
    end

    reg [7:0] out2816;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2816 = in0;
    end

    reg [7:0] out2817;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2817 = in0;
    end

    reg [7:0] out2818;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2818 = in0;
    end

    reg [7:0] out2819;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2819 = in0;
    end

    reg [7:0] out2820;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2820 = in0;
    end

    reg [7:0] out2821;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2821 = in0;
    end

    reg [7:0] out2822;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2822 = in0;
    end

    reg [7:0] out2823;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2823 = in0;
    end

    reg [7:0] out2824;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2824 = in0;
    end

    reg [7:0] out2825;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2825 = in0;
    end

    reg [7:0] out2826;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2826 = in0;
    end

    reg [7:0] out2827;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2827 = in0;
    end

    reg [7:0] out2828;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2828 = in0;
    end

    reg [7:0] out2829;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2829 = in0;
    end

    reg [7:0] out2830;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2830 = in0;
    end

    reg [7:0] out2831;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2831 = in0;
    end

    reg [7:0] out2832;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2832 = in0;
    end

    reg [7:0] out2833;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2833 = in0;
    end

    reg [7:0] out2834;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2834 = in0;
    end

    reg [7:0] out2835;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2835 = in0;
    end

    reg [7:0] out2836;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2836 = in0;
    end

    reg [7:0] out2837;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2837 = in0;
    end

    reg [7:0] out2838;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2838 = in0;
    end

    reg [7:0] out2839;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2839 = in0;
    end

    reg [7:0] out2840;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2840 = in0;
    end

    reg [7:0] out2841;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2841 = in0;
    end

    reg [7:0] out2842;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2842 = in0;
    end

    reg [7:0] out2843;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2843 = in0;
    end

    reg [7:0] out2844;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2844 = in0;
    end

    reg [7:0] out2845;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2845 = in0;
    end

    reg [7:0] out2846;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2846 = in0;
    end

    reg [7:0] out2847;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2847 = in0;
    end

    reg [7:0] out2848;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2848 = in0;
    end

    reg [7:0] out2849;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2849 = in0;
    end

    reg [7:0] out2850;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2850 = in0;
    end

    reg [7:0] out2851;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2851 = in0;
    end

    reg [7:0] out2852;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2852 = in0;
    end

    reg [7:0] out2853;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2853 = in0;
    end

    reg [7:0] out2854;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2854 = in0;
    end

    reg [7:0] out2855;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2855 = in0;
    end

    reg [7:0] out2856;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2856 = in0;
    end

    reg [7:0] out2857;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2857 = in0;
    end

    reg [7:0] out2858;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2858 = in0;
    end

    reg [7:0] out2859;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2859 = in0;
    end

    reg [7:0] out2860;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2860 = in0;
    end

    reg [7:0] out2861;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2861 = in0;
    end

    reg [7:0] out2862;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2862 = in0;
    end

    reg [7:0] out2863;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2863 = in0;
    end

    reg [7:0] out2864;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2864 = in0;
    end

    reg [7:0] out2865;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2865 = in0;
    end

    reg [7:0] out2866;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2866 = in0;
    end

    reg [7:0] out2867;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2867 = in0;
    end

    reg [7:0] out2868;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2868 = in0;
    end

    reg [7:0] out2869;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2869 = in0;
    end

    reg [7:0] out2870;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2870 = in0;
    end

    reg [7:0] out2871;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2871 = in0;
    end

    reg [7:0] out2872;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2872 = in0;
    end

    reg [7:0] out2873;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2873 = in0;
    end

    reg [7:0] out2874;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2874 = in0;
    end

    reg [7:0] out2875;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2875 = in0;
    end

    reg [7:0] out2876;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2876 = in0;
    end

    reg [7:0] out2877;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2877 = in0;
    end

    reg [7:0] out2878;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2878 = in0;
    end

    reg [7:0] out2879;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2879 = in0;
    end

    reg [7:0] out2880;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2880 = in0;
    end

    reg [7:0] out2881;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2881 = in0;
    end

    reg [7:0] out2882;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2882 = in0;
    end

    reg [7:0] out2883;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2883 = in0;
    end

    reg [7:0] out2884;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2884 = in0;
    end

    reg [7:0] out2885;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2885 = in0;
    end

    reg [7:0] out2886;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2886 = in0;
    end

    reg [7:0] out2887;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2887 = in0;
    end

    reg [7:0] out2888;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2888 = in0;
    end

    reg [7:0] out2889;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2889 = in0;
    end

    reg [7:0] out2890;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2890 = in0;
    end

    reg [7:0] out2891;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2891 = in0;
    end

    reg [7:0] out2892;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2892 = in0;
    end

    reg [7:0] out2893;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2893 = in0;
    end

    reg [7:0] out2894;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2894 = in0;
    end

    reg [7:0] out2895;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2895 = in0;
    end

    reg [7:0] out2896;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2896 = in0;
    end

    reg [7:0] out2897;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2897 = in0;
    end

    reg [7:0] out2898;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2898 = in0;
    end

    reg [7:0] out2899;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2899 = in0;
    end

    reg [7:0] out2900;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2900 = in0;
    end

    reg [7:0] out2901;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2901 = in0;
    end

    reg [7:0] out2902;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2902 = in0;
    end

    reg [7:0] out2903;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2903 = in0;
    end

    reg [7:0] out2904;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2904 = in0;
    end

    reg [7:0] out2905;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2905 = in0;
    end

    reg [7:0] out2906;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2906 = in0;
    end

    reg [7:0] out2907;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2907 = in0;
    end

    reg [7:0] out2908;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2908 = in0;
    end

    reg [7:0] out2909;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2909 = in0;
    end

    reg [7:0] out2910;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2910 = in0;
    end

    reg [7:0] out2911;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2911 = in0;
    end

    reg [7:0] out2912;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2912 = in0;
    end

    reg [7:0] out2913;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2913 = in0;
    end

    reg [7:0] out2914;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2914 = in0;
    end

    reg [7:0] out2915;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2915 = in0;
    end

    reg [7:0] out2916;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2916 = in0;
    end

    reg [7:0] out2917;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2917 = in0;
    end

    reg [7:0] out2918;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2918 = in0;
    end

    reg [7:0] out2919;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2919 = in0;
    end

    reg [7:0] out2920;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2920 = in0;
    end

    reg [7:0] out2921;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2921 = in0;
    end

    reg [7:0] out2922;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2922 = in0;
    end

    reg [7:0] out2923;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2923 = in0;
    end

    reg [7:0] out2924;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2924 = in0;
    end

    reg [7:0] out2925;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2925 = in0;
    end

    reg [7:0] out2926;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2926 = in0;
    end

    reg [7:0] out2927;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2927 = in0;
    end

    reg [7:0] out2928;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2928 = in0;
    end

    reg [7:0] out2929;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2929 = in0;
    end

    reg [7:0] out2930;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2930 = in0;
    end

    reg [7:0] out2931;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2931 = in0;
    end

    reg [7:0] out2932;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2932 = in0;
    end

    reg [7:0] out2933;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2933 = in0;
    end

    reg [7:0] out2934;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2934 = in0;
    end

    reg [7:0] out2935;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2935 = in0;
    end

    reg [7:0] out2936;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2936 = in0;
    end

    reg [7:0] out2937;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2937 = in0;
    end

    reg [7:0] out2938;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2938 = in0;
    end

    reg [7:0] out2939;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2939 = in0;
    end

    reg [7:0] out2940;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2940 = in0;
    end

    reg [7:0] out2941;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2941 = in0;
    end

    reg [7:0] out2942;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2942 = in0;
    end

    reg [7:0] out2943;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2943 = in0;
    end

    reg [7:0] out2944;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2944 = in0;
    end

    reg [7:0] out2945;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2945 = in0;
    end

    reg [7:0] out2946;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2946 = in0;
    end

    reg [7:0] out2947;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2947 = in0;
    end

    reg [7:0] out2948;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2948 = in0;
    end

    reg [7:0] out2949;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2949 = in0;
    end

    reg [7:0] out2950;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2950 = in0;
    end

    reg [7:0] out2951;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2951 = in0;
    end

    reg [7:0] out2952;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2952 = in0;
    end

    reg [7:0] out2953;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2953 = in0;
    end

    reg [7:0] out2954;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2954 = in0;
    end

    reg [7:0] out2955;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2955 = in0;
    end

    reg [7:0] out2956;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2956 = in0;
    end

    reg [7:0] out2957;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2957 = in0;
    end

    reg [7:0] out2958;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2958 = in0;
    end

    reg [7:0] out2959;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2959 = in0;
    end

    reg [7:0] out2960;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2960 = in0;
    end

    reg [7:0] out2961;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2961 = in0;
    end

    reg [7:0] out2962;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2962 = in0;
    end

    reg [7:0] out2963;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2963 = in0;
    end

    reg [7:0] out2964;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2964 = in0;
    end

    reg [7:0] out2965;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2965 = in0;
    end

    reg [7:0] out2966;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2966 = in0;
    end

    reg [7:0] out2967;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2967 = in0;
    end

    reg [7:0] out2968;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2968 = in0;
    end

    reg [7:0] out2969;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2969 = in0;
    end

    reg [7:0] out2970;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2970 = in0;
    end

    reg [7:0] out2971;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2971 = in0;
    end

    reg [7:0] out2972;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2972 = in0;
    end

    reg [7:0] out2973;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2973 = in0;
    end

    reg [7:0] out2974;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2974 = in0;
    end

    reg [7:0] out2975;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2975 = in0;
    end

    reg [7:0] out2976;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2976 = in0;
    end

    reg [7:0] out2977;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2977 = in0;
    end

    reg [7:0] out2978;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2978 = in0;
    end

    reg [7:0] out2979;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2979 = in0;
    end

    reg [7:0] out2980;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2980 = in0;
    end

    reg [7:0] out2981;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2981 = in0;
    end

    reg [7:0] out2982;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2982 = in0;
    end

    reg [7:0] out2983;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2983 = in0;
    end

    reg [7:0] out2984;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2984 = in0;
    end

    reg [7:0] out2985;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2985 = in0;
    end

    reg [7:0] out2986;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2986 = in0;
    end

    reg [7:0] out2987;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2987 = in0;
    end

    reg [7:0] out2988;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2988 = in0;
    end

    reg [7:0] out2989;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2989 = in0;
    end

    reg [7:0] out2990;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2990 = in0;
    end

    reg [7:0] out2991;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2991 = in0;
    end

    reg [7:0] out2992;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2992 = in0;
    end

    reg [7:0] out2993;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2993 = in0;
    end

    reg [7:0] out2994;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2994 = in0;
    end

    reg [7:0] out2995;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2995 = in0;
    end

    reg [7:0] out2996;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2996 = in0;
    end

    reg [7:0] out2997;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2997 = in0;
    end

    reg [7:0] out2998;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2998 = in0;
    end

    reg [7:0] out2999;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out2999 = in0;
    end

    reg [7:0] out3000;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3000 = in0;
    end

    reg [7:0] out3001;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3001 = in0;
    end

    reg [7:0] out3002;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3002 = in0;
    end

    reg [7:0] out3003;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3003 = in0;
    end

    reg [7:0] out3004;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3004 = in0;
    end

    reg [7:0] out3005;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3005 = in0;
    end

    reg [7:0] out3006;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3006 = in0;
    end

    reg [7:0] out3007;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3007 = in0;
    end

    reg [7:0] out3008;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3008 = in0;
    end

    reg [7:0] out3009;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3009 = in0;
    end

    reg [7:0] out3010;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3010 = in0;
    end

    reg [7:0] out3011;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3011 = in0;
    end

    reg [7:0] out3012;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3012 = in0;
    end

    reg [7:0] out3013;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3013 = in0;
    end

    reg [7:0] out3014;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3014 = in0;
    end

    reg [7:0] out3015;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3015 = in0;
    end

    reg [7:0] out3016;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3016 = in0;
    end

    reg [7:0] out3017;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3017 = in0;
    end

    reg [7:0] out3018;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3018 = in0;
    end

    reg [7:0] out3019;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3019 = in0;
    end

    reg [7:0] out3020;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3020 = in0;
    end

    reg [7:0] out3021;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3021 = in0;
    end

    reg [7:0] out3022;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3022 = in0;
    end

    reg [7:0] out3023;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3023 = in0;
    end

    reg [7:0] out3024;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3024 = in0;
    end

    reg [7:0] out3025;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3025 = in0;
    end

    reg [7:0] out3026;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3026 = in0;
    end

    reg [7:0] out3027;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3027 = in0;
    end

    reg [7:0] out3028;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3028 = in0;
    end

    reg [7:0] out3029;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3029 = in0;
    end

    reg [7:0] out3030;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3030 = in0;
    end

    reg [7:0] out3031;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3031 = in0;
    end

    reg [7:0] out3032;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3032 = in0;
    end

    reg [7:0] out3033;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3033 = in0;
    end

    reg [7:0] out3034;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3034 = in0;
    end

    reg [7:0] out3035;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3035 = in0;
    end

    reg [7:0] out3036;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3036 = in0;
    end

    reg [7:0] out3037;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3037 = in0;
    end

    reg [7:0] out3038;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3038 = in0;
    end

    reg [7:0] out3039;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3039 = in0;
    end

    reg [7:0] out3040;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3040 = in0;
    end

    reg [7:0] out3041;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3041 = in0;
    end

    reg [7:0] out3042;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3042 = in0;
    end

    reg [7:0] out3043;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3043 = in0;
    end

    reg [7:0] out3044;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3044 = in0;
    end

    reg [7:0] out3045;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3045 = in0;
    end

    reg [7:0] out3046;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3046 = in0;
    end

    reg [7:0] out3047;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3047 = in0;
    end

    reg [7:0] out3048;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3048 = in0;
    end

    reg [7:0] out3049;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3049 = in0;
    end

    reg [7:0] out3050;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3050 = in0;
    end

    reg [7:0] out3051;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3051 = in0;
    end

    reg [7:0] out3052;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3052 = in0;
    end

    reg [7:0] out3053;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3053 = in0;
    end

    reg [7:0] out3054;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3054 = in0;
    end

    reg [7:0] out3055;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3055 = in0;
    end

    reg [7:0] out3056;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3056 = in0;
    end

    reg [7:0] out3057;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3057 = in0;
    end

    reg [7:0] out3058;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3058 = in0;
    end

    reg [7:0] out3059;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3059 = in0;
    end

    reg [7:0] out3060;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3060 = in0;
    end

    reg [7:0] out3061;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3061 = in0;
    end

    reg [7:0] out3062;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3062 = in0;
    end

    reg [7:0] out3063;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3063 = in0;
    end

    reg [7:0] out3064;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3064 = in0;
    end

    reg [7:0] out3065;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3065 = in0;
    end

    reg [7:0] out3066;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3066 = in0;
    end

    reg [7:0] out3067;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3067 = in0;
    end

    reg [7:0] out3068;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3068 = in0;
    end

    reg [7:0] out3069;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3069 = in0;
    end

    reg [7:0] out3070;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3070 = in0;
    end

    reg [7:0] out3071;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3071 = in0;
    end

    reg [7:0] out3072;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3072 = in0;
    end

    reg [7:0] out3073;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3073 = in0;
    end

    reg [7:0] out3074;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3074 = in0;
    end

    reg [7:0] out3075;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3075 = in0;
    end

    reg [7:0] out3076;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3076 = in0;
    end

    reg [7:0] out3077;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3077 = in0;
    end

    reg [7:0] out3078;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3078 = in0;
    end

    reg [7:0] out3079;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3079 = in0;
    end

    reg [7:0] out3080;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3080 = in0;
    end

    reg [7:0] out3081;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3081 = in0;
    end

    reg [7:0] out3082;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3082 = in0;
    end

    reg [7:0] out3083;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3083 = in0;
    end

    reg [7:0] out3084;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3084 = in0;
    end

    reg [7:0] out3085;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3085 = in0;
    end

    reg [7:0] out3086;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3086 = in0;
    end

    reg [7:0] out3087;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3087 = in0;
    end

    reg [7:0] out3088;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3088 = in0;
    end

    reg [7:0] out3089;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3089 = in0;
    end

    reg [7:0] out3090;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3090 = in0;
    end

    reg [7:0] out3091;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3091 = in0;
    end

    reg [7:0] out3092;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3092 = in0;
    end

    reg [7:0] out3093;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3093 = in0;
    end

    reg [7:0] out3094;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3094 = in0;
    end

    reg [7:0] out3095;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3095 = in0;
    end

    reg [7:0] out3096;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3096 = in0;
    end

    reg [7:0] out3097;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3097 = in0;
    end

    reg [7:0] out3098;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3098 = in0;
    end

    reg [7:0] out3099;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3099 = in0;
    end

    reg [7:0] out3100;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3100 = in0;
    end

    reg [7:0] out3101;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3101 = in0;
    end

    reg [7:0] out3102;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3102 = in0;
    end

    reg [7:0] out3103;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3103 = in0;
    end

    reg [7:0] out3104;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3104 = in0;
    end

    reg [7:0] out3105;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3105 = in0;
    end

    reg [7:0] out3106;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3106 = in0;
    end

    reg [7:0] out3107;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3107 = in0;
    end

    reg [7:0] out3108;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3108 = in0;
    end

    reg [7:0] out3109;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3109 = in0;
    end

    reg [7:0] out3110;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3110 = in0;
    end

    reg [7:0] out3111;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3111 = in0;
    end

    reg [7:0] out3112;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3112 = in0;
    end

    reg [7:0] out3113;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3113 = in0;
    end

    reg [7:0] out3114;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3114 = in0;
    end

    reg [7:0] out3115;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3115 = in0;
    end

    reg [7:0] out3116;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3116 = in0;
    end

    reg [7:0] out3117;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3117 = in0;
    end

    reg [7:0] out3118;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3118 = in0;
    end

    reg [7:0] out3119;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3119 = in0;
    end

    reg [7:0] out3120;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3120 = in0;
    end

    reg [7:0] out3121;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3121 = in0;
    end

    reg [7:0] out3122;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3122 = in0;
    end

    reg [7:0] out3123;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3123 = in0;
    end

    reg [7:0] out3124;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3124 = in0;
    end

    reg [7:0] out3125;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3125 = in0;
    end

    reg [7:0] out3126;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3126 = in0;
    end

    reg [7:0] out3127;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3127 = in0;
    end

    reg [7:0] out3128;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3128 = in0;
    end

    reg [7:0] out3129;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3129 = in0;
    end

    reg [7:0] out3130;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3130 = in0;
    end

    reg [7:0] out3131;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3131 = in0;
    end

    reg [7:0] out3132;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3132 = in0;
    end

    reg [7:0] out3133;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3133 = in0;
    end

    reg [7:0] out3134;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3134 = in0;
    end

    reg [7:0] out3135;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3135 = in0;
    end

    reg [7:0] out3136;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3136 = in0;
    end

    reg [7:0] out3137;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3137 = in0;
    end

    reg [7:0] out3138;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3138 = in0;
    end

    reg [7:0] out3139;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3139 = in0;
    end

    reg [7:0] out3140;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3140 = in0;
    end

    reg [7:0] out3141;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3141 = in0;
    end

    reg [7:0] out3142;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3142 = in0;
    end

    reg [7:0] out3143;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3143 = in0;
    end

    reg [7:0] out3144;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3144 = in0;
    end

    reg [7:0] out3145;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3145 = in0;
    end

    reg [7:0] out3146;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3146 = in0;
    end

    reg [7:0] out3147;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3147 = in0;
    end

    reg [7:0] out3148;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3148 = in0;
    end

    reg [7:0] out3149;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3149 = in0;
    end

    reg [7:0] out3150;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3150 = in0;
    end

    reg [7:0] out3151;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3151 = in0;
    end

    reg [7:0] out3152;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3152 = in0;
    end

    reg [7:0] out3153;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3153 = in0;
    end

    reg [7:0] out3154;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3154 = in0;
    end

    reg [7:0] out3155;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3155 = in0;
    end

    reg [7:0] out3156;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3156 = in0;
    end

    reg [7:0] out3157;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3157 = in0;
    end

    reg [7:0] out3158;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3158 = in0;
    end

    reg [7:0] out3159;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3159 = in0;
    end

    reg [7:0] out3160;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3160 = in0;
    end

    reg [7:0] out3161;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3161 = in0;
    end

    reg [7:0] out3162;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3162 = in0;
    end

    reg [7:0] out3163;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3163 = in0;
    end

    reg [7:0] out3164;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3164 = in0;
    end

    reg [7:0] out3165;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3165 = in0;
    end

    reg [7:0] out3166;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3166 = in0;
    end

    reg [7:0] out3167;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3167 = in0;
    end

    reg [7:0] out3168;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3168 = in0;
    end

    reg [7:0] out3169;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3169 = in0;
    end

    reg [7:0] out3170;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3170 = in0;
    end

    reg [7:0] out3171;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3171 = in0;
    end

    reg [7:0] out3172;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3172 = in0;
    end

    reg [7:0] out3173;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3173 = in0;
    end

    reg [7:0] out3174;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3174 = in0;
    end

    reg [7:0] out3175;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3175 = in0;
    end

    reg [7:0] out3176;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3176 = in0;
    end

    reg [7:0] out3177;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3177 = in0;
    end

    reg [7:0] out3178;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3178 = in0;
    end

    reg [7:0] out3179;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3179 = in0;
    end

    reg [7:0] out3180;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3180 = in0;
    end

    reg [7:0] out3181;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3181 = in0;
    end

    reg [7:0] out3182;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3182 = in0;
    end

    reg [7:0] out3183;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3183 = in0;
    end

    reg [7:0] out3184;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3184 = in0;
    end

    reg [7:0] out3185;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3185 = in0;
    end

    reg [7:0] out3186;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3186 = in0;
    end

    reg [7:0] out3187;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3187 = in0;
    end

    reg [7:0] out3188;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3188 = in0;
    end

    reg [7:0] out3189;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3189 = in0;
    end

    reg [7:0] out3190;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3190 = in0;
    end

    reg [7:0] out3191;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3191 = in0;
    end

    reg [7:0] out3192;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3192 = in0;
    end

    reg [7:0] out3193;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3193 = in0;
    end

    reg [7:0] out3194;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3194 = in0;
    end

    reg [7:0] out3195;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3195 = in0;
    end

    reg [7:0] out3196;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3196 = in0;
    end

    reg [7:0] out3197;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3197 = in0;
    end

    reg [7:0] out3198;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3198 = in0;
    end

    reg [7:0] out3199;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3199 = in0;
    end

    reg [7:0] out3200;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3200 = in0;
    end

    reg [7:0] out3201;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3201 = in0;
    end

    reg [7:0] out3202;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3202 = in0;
    end

    reg [7:0] out3203;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3203 = in0;
    end

    reg [7:0] out3204;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3204 = in0;
    end

    reg [7:0] out3205;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3205 = in0;
    end

    reg [7:0] out3206;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3206 = in0;
    end

    reg [7:0] out3207;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3207 = in0;
    end

    reg [7:0] out3208;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3208 = in0;
    end

    reg [7:0] out3209;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3209 = in0;
    end

    reg [7:0] out3210;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3210 = in0;
    end

    reg [7:0] out3211;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3211 = in0;
    end

    reg [7:0] out3212;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3212 = in0;
    end

    reg [7:0] out3213;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3213 = in0;
    end

    reg [7:0] out3214;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3214 = in0;
    end

    reg [7:0] out3215;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3215 = in0;
    end

    reg [7:0] out3216;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3216 = in0;
    end

    reg [7:0] out3217;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3217 = in0;
    end

    reg [7:0] out3218;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3218 = in0;
    end

    reg [7:0] out3219;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3219 = in0;
    end

    reg [7:0] out3220;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3220 = in0;
    end

    reg [7:0] out3221;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3221 = in0;
    end

    reg [7:0] out3222;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3222 = in0;
    end

    reg [7:0] out3223;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3223 = in0;
    end

    reg [7:0] out3224;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3224 = in0;
    end

    reg [7:0] out3225;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3225 = in0;
    end

    reg [7:0] out3226;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3226 = in0;
    end

    reg [7:0] out3227;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3227 = in0;
    end

    reg [7:0] out3228;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3228 = in0;
    end

    reg [7:0] out3229;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3229 = in0;
    end

    reg [7:0] out3230;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3230 = in0;
    end

    reg [7:0] out3231;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3231 = in0;
    end

    reg [7:0] out3232;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3232 = in0;
    end

    reg [7:0] out3233;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3233 = in0;
    end

    reg [7:0] out3234;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3234 = in0;
    end

    reg [7:0] out3235;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3235 = in0;
    end

    reg [7:0] out3236;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3236 = in0;
    end

    reg [7:0] out3237;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3237 = in0;
    end

    reg [7:0] out3238;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3238 = in0;
    end

    reg [7:0] out3239;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3239 = in0;
    end

    reg [7:0] out3240;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3240 = in0;
    end

    reg [7:0] out3241;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3241 = in0;
    end

    reg [7:0] out3242;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3242 = in0;
    end

    reg [7:0] out3243;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3243 = in0;
    end

    reg [7:0] out3244;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3244 = in0;
    end

    reg [7:0] out3245;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3245 = in0;
    end

    reg [7:0] out3246;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3246 = in0;
    end

    reg [7:0] out3247;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3247 = in0;
    end

    reg [7:0] out3248;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3248 = in0;
    end

    reg [7:0] out3249;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3249 = in0;
    end

    reg [7:0] out3250;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3250 = in0;
    end

    reg [7:0] out3251;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3251 = in0;
    end

    reg [7:0] out3252;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3252 = in0;
    end

    reg [7:0] out3253;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3253 = in0;
    end

    reg [7:0] out3254;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3254 = in0;
    end

    reg [7:0] out3255;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3255 = in0;
    end

    reg [7:0] out3256;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3256 = in0;
    end

    reg [7:0] out3257;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3257 = in0;
    end

    reg [7:0] out3258;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3258 = in0;
    end

    reg [7:0] out3259;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3259 = in0;
    end

    reg [7:0] out3260;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3260 = in0;
    end

    reg [7:0] out3261;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3261 = in0;
    end

    reg [7:0] out3262;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3262 = in0;
    end

    reg [7:0] out3263;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3263 = in0;
    end

    reg [7:0] out3264;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3264 = in0;
    end

    reg [7:0] out3265;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3265 = in0;
    end

    reg [7:0] out3266;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3266 = in0;
    end

    reg [7:0] out3267;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3267 = in0;
    end

    reg [7:0] out3268;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3268 = in0;
    end

    reg [7:0] out3269;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3269 = in0;
    end

    reg [7:0] out3270;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3270 = in0;
    end

    reg [7:0] out3271;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3271 = in0;
    end

    reg [7:0] out3272;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3272 = in0;
    end

    reg [7:0] out3273;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3273 = in0;
    end

    reg [7:0] out3274;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3274 = in0;
    end

    reg [7:0] out3275;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3275 = in0;
    end

    reg [7:0] out3276;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3276 = in0;
    end

    reg [7:0] out3277;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3277 = in0;
    end

    reg [7:0] out3278;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3278 = in0;
    end

    reg [7:0] out3279;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3279 = in0;
    end

    reg [7:0] out3280;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3280 = in0;
    end

    reg [7:0] out3281;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3281 = in0;
    end

    reg [7:0] out3282;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3282 = in0;
    end

    reg [7:0] out3283;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3283 = in0;
    end

    reg [7:0] out3284;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3284 = in0;
    end

    reg [7:0] out3285;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3285 = in0;
    end

    reg [7:0] out3286;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3286 = in0;
    end

    reg [7:0] out3287;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3287 = in0;
    end

    reg [7:0] out3288;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3288 = in0;
    end

    reg [7:0] out3289;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3289 = in0;
    end

    reg [7:0] out3290;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3290 = in0;
    end

    reg [7:0] out3291;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3291 = in0;
    end

    reg [7:0] out3292;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3292 = in0;
    end

    reg [7:0] out3293;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3293 = in0;
    end

    reg [7:0] out3294;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3294 = in0;
    end

    reg [7:0] out3295;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3295 = in0;
    end

    reg [7:0] out3296;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3296 = in0;
    end

    reg [7:0] out3297;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3297 = in0;
    end

    reg [7:0] out3298;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3298 = in0;
    end

    reg [7:0] out3299;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3299 = in0;
    end

    reg [7:0] out3300;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3300 = in0;
    end

    reg [7:0] out3301;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3301 = in0;
    end

    reg [7:0] out3302;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3302 = in0;
    end

    reg [7:0] out3303;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3303 = in0;
    end

    reg [7:0] out3304;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3304 = in0;
    end

    reg [7:0] out3305;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3305 = in0;
    end

    reg [7:0] out3306;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3306 = in0;
    end

    reg [7:0] out3307;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3307 = in0;
    end

    reg [7:0] out3308;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3308 = in0;
    end

    reg [7:0] out3309;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3309 = in0;
    end

    reg [7:0] out3310;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3310 = in0;
    end

    reg [7:0] out3311;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3311 = in0;
    end

    reg [7:0] out3312;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3312 = in0;
    end

    reg [7:0] out3313;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3313 = in0;
    end

    reg [7:0] out3314;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3314 = in0;
    end

    reg [7:0] out3315;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3315 = in0;
    end

    reg [7:0] out3316;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3316 = in0;
    end

    reg [7:0] out3317;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3317 = in0;
    end

    reg [7:0] out3318;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3318 = in0;
    end

    reg [7:0] out3319;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3319 = in0;
    end

    reg [7:0] out3320;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3320 = in0;
    end

    reg [7:0] out3321;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3321 = in0;
    end

    reg [7:0] out3322;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3322 = in0;
    end

    reg [7:0] out3323;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3323 = in0;
    end

    reg [7:0] out3324;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3324 = in0;
    end

    reg [7:0] out3325;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3325 = in0;
    end

    reg [7:0] out3326;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3326 = in0;
    end

    reg [7:0] out3327;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3327 = in0;
    end

    reg [7:0] out3328;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3328 = in0;
    end

    reg [7:0] out3329;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3329 = in0;
    end

    reg [7:0] out3330;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3330 = in0;
    end

    reg [7:0] out3331;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3331 = in0;
    end

    reg [7:0] out3332;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3332 = in0;
    end

    reg [7:0] out3333;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3333 = in0;
    end

    reg [7:0] out3334;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3334 = in0;
    end

    reg [7:0] out3335;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3335 = in0;
    end

    reg [7:0] out3336;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3336 = in0;
    end

    reg [7:0] out3337;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3337 = in0;
    end

    reg [7:0] out3338;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3338 = in0;
    end

    reg [7:0] out3339;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3339 = in0;
    end

    reg [7:0] out3340;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3340 = in0;
    end

    reg [7:0] out3341;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3341 = in0;
    end

    reg [7:0] out3342;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3342 = in0;
    end

    reg [7:0] out3343;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3343 = in0;
    end

    reg [7:0] out3344;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3344 = in0;
    end

    reg [7:0] out3345;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3345 = in0;
    end

    reg [7:0] out3346;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3346 = in0;
    end

    reg [7:0] out3347;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3347 = in0;
    end

    reg [7:0] out3348;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3348 = in0;
    end

    reg [7:0] out3349;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3349 = in0;
    end

    reg [7:0] out3350;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3350 = in0;
    end

    reg [7:0] out3351;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3351 = in0;
    end

    reg [7:0] out3352;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3352 = in0;
    end

    reg [7:0] out3353;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3353 = in0;
    end

    reg [7:0] out3354;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3354 = in0;
    end

    reg [7:0] out3355;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3355 = in0;
    end

    reg [7:0] out3356;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3356 = in0;
    end

    reg [7:0] out3357;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3357 = in0;
    end

    reg [7:0] out3358;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3358 = in0;
    end

    reg [7:0] out3359;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3359 = in0;
    end

    reg [7:0] out3360;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3360 = in0;
    end

    reg [7:0] out3361;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3361 = in0;
    end

    reg [7:0] out3362;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3362 = in0;
    end

    reg [7:0] out3363;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3363 = in0;
    end

    reg [7:0] out3364;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3364 = in0;
    end

    reg [7:0] out3365;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3365 = in0;
    end

    reg [7:0] out3366;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3366 = in0;
    end

    reg [7:0] out3367;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3367 = in0;
    end

    reg [7:0] out3368;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3368 = in0;
    end

    reg [7:0] out3369;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3369 = in0;
    end

    reg [7:0] out3370;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3370 = in0;
    end

    reg [7:0] out3371;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3371 = in0;
    end

    reg [7:0] out3372;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3372 = in0;
    end

    reg [7:0] out3373;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3373 = in0;
    end

    reg [7:0] out3374;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3374 = in0;
    end

    reg [7:0] out3375;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3375 = in0;
    end

    reg [7:0] out3376;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3376 = in0;
    end

    reg [7:0] out3377;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3377 = in0;
    end

    reg [7:0] out3378;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3378 = in0;
    end

    reg [7:0] out3379;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3379 = in0;
    end

    reg [7:0] out3380;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3380 = in0;
    end

    reg [7:0] out3381;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3381 = in0;
    end

    reg [7:0] out3382;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3382 = in0;
    end

    reg [7:0] out3383;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3383 = in0;
    end

    reg [7:0] out3384;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3384 = in0;
    end

    reg [7:0] out3385;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3385 = in0;
    end

    reg [7:0] out3386;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3386 = in0;
    end

    reg [7:0] out3387;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3387 = in0;
    end

    reg [7:0] out3388;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3388 = in0;
    end

    reg [7:0] out3389;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3389 = in0;
    end

    reg [7:0] out3390;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3390 = in0;
    end

    reg [7:0] out3391;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3391 = in0;
    end

    reg [7:0] out3392;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3392 = in0;
    end

    reg [7:0] out3393;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3393 = in0;
    end

    reg [7:0] out3394;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3394 = in0;
    end

    reg [7:0] out3395;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3395 = in0;
    end

    reg [7:0] out3396;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3396 = in0;
    end

    reg [7:0] out3397;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3397 = in0;
    end

    reg [7:0] out3398;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3398 = in0;
    end

    reg [7:0] out3399;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3399 = in0;
    end

    reg [7:0] out3400;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3400 = in0;
    end

    reg [7:0] out3401;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3401 = in0;
    end

    reg [7:0] out3402;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3402 = in0;
    end

    reg [7:0] out3403;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3403 = in0;
    end

    reg [7:0] out3404;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3404 = in0;
    end

    reg [7:0] out3405;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3405 = in0;
    end

    reg [7:0] out3406;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3406 = in0;
    end

    reg [7:0] out3407;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3407 = in0;
    end

    reg [7:0] out3408;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3408 = in0;
    end

    reg [7:0] out3409;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3409 = in0;
    end

    reg [7:0] out3410;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3410 = in0;
    end

    reg [7:0] out3411;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3411 = in0;
    end

    reg [7:0] out3412;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3412 = in0;
    end

    reg [7:0] out3413;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3413 = in0;
    end

    reg [7:0] out3414;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3414 = in0;
    end

    reg [7:0] out3415;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3415 = in0;
    end

    reg [7:0] out3416;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3416 = in0;
    end

    reg [7:0] out3417;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3417 = in0;
    end

    reg [7:0] out3418;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3418 = in0;
    end

    reg [7:0] out3419;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3419 = in0;
    end

    reg [7:0] out3420;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3420 = in0;
    end

    reg [7:0] out3421;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3421 = in0;
    end

    reg [7:0] out3422;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3422 = in0;
    end

    reg [7:0] out3423;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3423 = in0;
    end

    reg [7:0] out3424;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3424 = in0;
    end

    reg [7:0] out3425;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3425 = in0;
    end

    reg [7:0] out3426;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3426 = in0;
    end

    reg [7:0] out3427;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3427 = in0;
    end

    reg [7:0] out3428;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3428 = in0;
    end

    reg [7:0] out3429;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3429 = in0;
    end

    reg [7:0] out3430;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3430 = in0;
    end

    reg [7:0] out3431;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3431 = in0;
    end

    reg [7:0] out3432;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3432 = in0;
    end

    reg [7:0] out3433;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3433 = in0;
    end

    reg [7:0] out3434;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3434 = in0;
    end

    reg [7:0] out3435;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3435 = in0;
    end

    reg [7:0] out3436;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3436 = in0;
    end

    reg [7:0] out3437;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3437 = in0;
    end

    reg [7:0] out3438;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3438 = in0;
    end

    reg [7:0] out3439;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3439 = in0;
    end

    reg [7:0] out3440;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3440 = in0;
    end

    reg [7:0] out3441;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3441 = in0;
    end

    reg [7:0] out3442;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3442 = in0;
    end

    reg [7:0] out3443;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3443 = in0;
    end

    reg [7:0] out3444;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3444 = in0;
    end

    reg [7:0] out3445;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3445 = in0;
    end

    reg [7:0] out3446;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3446 = in0;
    end

    reg [7:0] out3447;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3447 = in0;
    end

    reg [7:0] out3448;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3448 = in0;
    end

    reg [7:0] out3449;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3449 = in0;
    end

    reg [7:0] out3450;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3450 = in0;
    end

    reg [7:0] out3451;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3451 = in0;
    end

    reg [7:0] out3452;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3452 = in0;
    end

    reg [7:0] out3453;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3453 = in0;
    end

    reg [7:0] out3454;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3454 = in0;
    end

    reg [7:0] out3455;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3455 = in0;
    end

    reg [7:0] out3456;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3456 = in0;
    end

    reg [7:0] out3457;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3457 = in0;
    end

    reg [7:0] out3458;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3458 = in0;
    end

    reg [7:0] out3459;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3459 = in0;
    end

    reg [7:0] out3460;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3460 = in0;
    end

    reg [7:0] out3461;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3461 = in0;
    end

    reg [7:0] out3462;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3462 = in0;
    end

    reg [7:0] out3463;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3463 = in0;
    end

    reg [7:0] out3464;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3464 = in0;
    end

    reg [7:0] out3465;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3465 = in0;
    end

    reg [7:0] out3466;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3466 = in0;
    end

    reg [7:0] out3467;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3467 = in0;
    end

    reg [7:0] out3468;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3468 = in0;
    end

    reg [7:0] out3469;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3469 = in0;
    end

    reg [7:0] out3470;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3470 = in0;
    end

    reg [7:0] out3471;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3471 = in0;
    end

    reg [7:0] out3472;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3472 = in0;
    end

    reg [7:0] out3473;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3473 = in0;
    end

    reg [7:0] out3474;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3474 = in0;
    end

    reg [7:0] out3475;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3475 = in0;
    end

    reg [7:0] out3476;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3476 = in0;
    end

    reg [7:0] out3477;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3477 = in0;
    end

    reg [7:0] out3478;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3478 = in0;
    end

    reg [7:0] out3479;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3479 = in0;
    end

    reg [7:0] out3480;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3480 = in0;
    end

    reg [7:0] out3481;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3481 = in0;
    end

    reg [7:0] out3482;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3482 = in0;
    end

    reg [7:0] out3483;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3483 = in0;
    end

    reg [7:0] out3484;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3484 = in0;
    end

    reg [7:0] out3485;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3485 = in0;
    end

    reg [7:0] out3486;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3486 = in0;
    end

    reg [7:0] out3487;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3487 = in0;
    end

    reg [7:0] out3488;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3488 = in0;
    end

    reg [7:0] out3489;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3489 = in0;
    end

    reg [7:0] out3490;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3490 = in0;
    end

    reg [7:0] out3491;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3491 = in0;
    end

    reg [7:0] out3492;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3492 = in0;
    end

    reg [7:0] out3493;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3493 = in0;
    end

    reg [7:0] out3494;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3494 = in0;
    end

    reg [7:0] out3495;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3495 = in0;
    end

    reg [7:0] out3496;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3496 = in0;
    end

    reg [7:0] out3497;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3497 = in0;
    end

    reg [7:0] out3498;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3498 = in0;
    end

    reg [7:0] out3499;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3499 = in0;
    end

    reg [7:0] out3500;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3500 = in0;
    end

    reg [7:0] out3501;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3501 = in0;
    end

    reg [7:0] out3502;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3502 = in0;
    end

    reg [7:0] out3503;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3503 = in0;
    end

    reg [7:0] out3504;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3504 = in0;
    end

    reg [7:0] out3505;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3505 = in0;
    end

    reg [7:0] out3506;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3506 = in0;
    end

    reg [7:0] out3507;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3507 = in0;
    end

    reg [7:0] out3508;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3508 = in0;
    end

    reg [7:0] out3509;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3509 = in0;
    end

    reg [7:0] out3510;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3510 = in0;
    end

    reg [7:0] out3511;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3511 = in0;
    end

    reg [7:0] out3512;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3512 = in0;
    end

    reg [7:0] out3513;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3513 = in0;
    end

    reg [7:0] out3514;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3514 = in0;
    end

    reg [7:0] out3515;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3515 = in0;
    end

    reg [7:0] out3516;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3516 = in0;
    end

    reg [7:0] out3517;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3517 = in0;
    end

    reg [7:0] out3518;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3518 = in0;
    end

    reg [7:0] out3519;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3519 = in0;
    end

    reg [7:0] out3520;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3520 = in0;
    end

    reg [7:0] out3521;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3521 = in0;
    end

    reg [7:0] out3522;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3522 = in0;
    end

    reg [7:0] out3523;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3523 = in0;
    end

    reg [7:0] out3524;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3524 = in0;
    end

    reg [7:0] out3525;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3525 = in0;
    end

    reg [7:0] out3526;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3526 = in0;
    end

    reg [7:0] out3527;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3527 = in0;
    end

    reg [7:0] out3528;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3528 = in0;
    end

    reg [7:0] out3529;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3529 = in0;
    end

    reg [7:0] out3530;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3530 = in0;
    end

    reg [7:0] out3531;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3531 = in0;
    end

    reg [7:0] out3532;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3532 = in0;
    end

    reg [7:0] out3533;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3533 = in0;
    end

    reg [7:0] out3534;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3534 = in0;
    end

    reg [7:0] out3535;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3535 = in0;
    end

    reg [7:0] out3536;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3536 = in0;
    end

    reg [7:0] out3537;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3537 = in0;
    end

    reg [7:0] out3538;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3538 = in0;
    end

    reg [7:0] out3539;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3539 = in0;
    end

    reg [7:0] out3540;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3540 = in0;
    end

    reg [7:0] out3541;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3541 = in0;
    end

    reg [7:0] out3542;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3542 = in0;
    end

    reg [7:0] out3543;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3543 = in0;
    end

    reg [7:0] out3544;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3544 = in0;
    end

    reg [7:0] out3545;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3545 = in0;
    end

    reg [7:0] out3546;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3546 = in0;
    end

    reg [7:0] out3547;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3547 = in0;
    end

    reg [7:0] out3548;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3548 = in0;
    end

    reg [7:0] out3549;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3549 = in0;
    end

    reg [7:0] out3550;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3550 = in0;
    end

    reg [7:0] out3551;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3551 = in0;
    end

    reg [7:0] out3552;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3552 = in0;
    end

    reg [7:0] out3553;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3553 = in0;
    end

    reg [7:0] out3554;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3554 = in0;
    end

    reg [7:0] out3555;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3555 = in0;
    end

    reg [7:0] out3556;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3556 = in0;
    end

    reg [7:0] out3557;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3557 = in0;
    end

    reg [7:0] out3558;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3558 = in0;
    end

    reg [7:0] out3559;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3559 = in0;
    end

    reg [7:0] out3560;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3560 = in0;
    end

    reg [7:0] out3561;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3561 = in0;
    end

    reg [7:0] out3562;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3562 = in0;
    end

    reg [7:0] out3563;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3563 = in0;
    end

    reg [7:0] out3564;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3564 = in0;
    end

    reg [7:0] out3565;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3565 = in0;
    end

    reg [7:0] out3566;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3566 = in0;
    end

    reg [7:0] out3567;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3567 = in0;
    end

    reg [7:0] out3568;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3568 = in0;
    end

    reg [7:0] out3569;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3569 = in0;
    end

    reg [7:0] out3570;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3570 = in0;
    end

    reg [7:0] out3571;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3571 = in0;
    end

    reg [7:0] out3572;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3572 = in0;
    end

    reg [7:0] out3573;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3573 = in0;
    end

    reg [7:0] out3574;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3574 = in0;
    end

    reg [7:0] out3575;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3575 = in0;
    end

    reg [7:0] out3576;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3576 = in0;
    end

    reg [7:0] out3577;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3577 = in0;
    end

    reg [7:0] out3578;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3578 = in0;
    end

    reg [7:0] out3579;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3579 = in0;
    end

    reg [7:0] out3580;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3580 = in0;
    end

    reg [7:0] out3581;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3581 = in0;
    end

    reg [7:0] out3582;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3582 = in0;
    end

    reg [7:0] out3583;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3583 = in0;
    end

    reg [7:0] out3584;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3584 = in0;
    end

    reg [7:0] out3585;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3585 = in0;
    end

    reg [7:0] out3586;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3586 = in0;
    end

    reg [7:0] out3587;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3587 = in0;
    end

    reg [7:0] out3588;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3588 = in0;
    end

    reg [7:0] out3589;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3589 = in0;
    end

    reg [7:0] out3590;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3590 = in0;
    end

    reg [7:0] out3591;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3591 = in0;
    end

    reg [7:0] out3592;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3592 = in0;
    end

    reg [7:0] out3593;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3593 = in0;
    end

    reg [7:0] out3594;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3594 = in0;
    end

    reg [7:0] out3595;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3595 = in0;
    end

    reg [7:0] out3596;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3596 = in0;
    end

    reg [7:0] out3597;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3597 = in0;
    end

    reg [7:0] out3598;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3598 = in0;
    end

    reg [7:0] out3599;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3599 = in0;
    end

    reg [7:0] out3600;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3600 = in0;
    end

    reg [7:0] out3601;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3601 = in0;
    end

    reg [7:0] out3602;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3602 = in0;
    end

    reg [7:0] out3603;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3603 = in0;
    end

    reg [7:0] out3604;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3604 = in0;
    end

    reg [7:0] out3605;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3605 = in0;
    end

    reg [7:0] out3606;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3606 = in0;
    end

    reg [7:0] out3607;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3607 = in0;
    end

    reg [7:0] out3608;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3608 = in0;
    end

    reg [7:0] out3609;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3609 = in0;
    end

    reg [7:0] out3610;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3610 = in0;
    end

    reg [7:0] out3611;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3611 = in0;
    end

    reg [7:0] out3612;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3612 = in0;
    end

    reg [7:0] out3613;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3613 = in0;
    end

    reg [7:0] out3614;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3614 = in0;
    end

    reg [7:0] out3615;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3615 = in0;
    end

    reg [7:0] out3616;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3616 = in0;
    end

    reg [7:0] out3617;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3617 = in0;
    end

    reg [7:0] out3618;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3618 = in0;
    end

    reg [7:0] out3619;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3619 = in0;
    end

    reg [7:0] out3620;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3620 = in0;
    end

    reg [7:0] out3621;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3621 = in0;
    end

    reg [7:0] out3622;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3622 = in0;
    end

    reg [7:0] out3623;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3623 = in0;
    end

    reg [7:0] out3624;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3624 = in0;
    end

    reg [7:0] out3625;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3625 = in0;
    end

    reg [7:0] out3626;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3626 = in0;
    end

    reg [7:0] out3627;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3627 = in0;
    end

    reg [7:0] out3628;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3628 = in0;
    end

    reg [7:0] out3629;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3629 = in0;
    end

    reg [7:0] out3630;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3630 = in0;
    end

    reg [7:0] out3631;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3631 = in0;
    end

    reg [7:0] out3632;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3632 = in0;
    end

    reg [7:0] out3633;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3633 = in0;
    end

    reg [7:0] out3634;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3634 = in0;
    end

    reg [7:0] out3635;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3635 = in0;
    end

    reg [7:0] out3636;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3636 = in0;
    end

    reg [7:0] out3637;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3637 = in0;
    end

    reg [7:0] out3638;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3638 = in0;
    end

    reg [7:0] out3639;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3639 = in0;
    end

    reg [7:0] out3640;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3640 = in0;
    end

    reg [7:0] out3641;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3641 = in0;
    end

    reg [7:0] out3642;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3642 = in0;
    end

    reg [7:0] out3643;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3643 = in0;
    end

    reg [7:0] out3644;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3644 = in0;
    end

    reg [7:0] out3645;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3645 = in0;
    end

    reg [7:0] out3646;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3646 = in0;
    end

    reg [7:0] out3647;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3647 = in0;
    end

    reg [7:0] out3648;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3648 = in0;
    end

    reg [7:0] out3649;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3649 = in0;
    end

    reg [7:0] out3650;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3650 = in0;
    end

    reg [7:0] out3651;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3651 = in0;
    end

    reg [7:0] out3652;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3652 = in0;
    end

    reg [7:0] out3653;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3653 = in0;
    end

    reg [7:0] out3654;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3654 = in0;
    end

    reg [7:0] out3655;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3655 = in0;
    end

    reg [7:0] out3656;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3656 = in0;
    end

    reg [7:0] out3657;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3657 = in0;
    end

    reg [7:0] out3658;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3658 = in0;
    end

    reg [7:0] out3659;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3659 = in0;
    end

    reg [7:0] out3660;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3660 = in0;
    end

    reg [7:0] out3661;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3661 = in0;
    end

    reg [7:0] out3662;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3662 = in0;
    end

    reg [7:0] out3663;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3663 = in0;
    end

    reg [7:0] out3664;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3664 = in0;
    end

    reg [7:0] out3665;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3665 = in0;
    end

    reg [7:0] out3666;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3666 = in0;
    end

    reg [7:0] out3667;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3667 = in0;
    end

    reg [7:0] out3668;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3668 = in0;
    end

    reg [7:0] out3669;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3669 = in0;
    end

    reg [7:0] out3670;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3670 = in0;
    end

    reg [7:0] out3671;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3671 = in0;
    end

    reg [7:0] out3672;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3672 = in0;
    end

    reg [7:0] out3673;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3673 = in0;
    end

    reg [7:0] out3674;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3674 = in0;
    end

    reg [7:0] out3675;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3675 = in0;
    end

    reg [7:0] out3676;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3676 = in0;
    end

    reg [7:0] out3677;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3677 = in0;
    end

    reg [7:0] out3678;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3678 = in0;
    end

    reg [7:0] out3679;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3679 = in0;
    end

    reg [7:0] out3680;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3680 = in0;
    end

    reg [7:0] out3681;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3681 = in0;
    end

    reg [7:0] out3682;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3682 = in0;
    end

    reg [7:0] out3683;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3683 = in0;
    end

    reg [7:0] out3684;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3684 = in0;
    end

    reg [7:0] out3685;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3685 = in0;
    end

    reg [7:0] out3686;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3686 = in0;
    end

    reg [7:0] out3687;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3687 = in0;
    end

    reg [7:0] out3688;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3688 = in0;
    end

    reg [7:0] out3689;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3689 = in0;
    end

    reg [7:0] out3690;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3690 = in0;
    end

    reg [7:0] out3691;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3691 = in0;
    end

    reg [7:0] out3692;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3692 = in0;
    end

    reg [7:0] out3693;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3693 = in0;
    end

    reg [7:0] out3694;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3694 = in0;
    end

    reg [7:0] out3695;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3695 = in0;
    end

    reg [7:0] out3696;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3696 = in0;
    end

    reg [7:0] out3697;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3697 = in0;
    end

    reg [7:0] out3698;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3698 = in0;
    end

    reg [7:0] out3699;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3699 = in0;
    end

    reg [7:0] out3700;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3700 = in0;
    end

    reg [7:0] out3701;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3701 = in0;
    end

    reg [7:0] out3702;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3702 = in0;
    end

    reg [7:0] out3703;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3703 = in0;
    end

    reg [7:0] out3704;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3704 = in0;
    end

    reg [7:0] out3705;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3705 = in0;
    end

    reg [7:0] out3706;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3706 = in0;
    end

    reg [7:0] out3707;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3707 = in0;
    end

    reg [7:0] out3708;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3708 = in0;
    end

    reg [7:0] out3709;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3709 = in0;
    end

    reg [7:0] out3710;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3710 = in0;
    end

    reg [7:0] out3711;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3711 = in0;
    end

    reg [7:0] out3712;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3712 = in0;
    end

    reg [7:0] out3713;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3713 = in0;
    end

    reg [7:0] out3714;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3714 = in0;
    end

    reg [7:0] out3715;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3715 = in0;
    end

    reg [7:0] out3716;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3716 = in0;
    end

    reg [7:0] out3717;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3717 = in0;
    end

    reg [7:0] out3718;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3718 = in0;
    end

    reg [7:0] out3719;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3719 = in0;
    end

    reg [7:0] out3720;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3720 = in0;
    end

    reg [7:0] out3721;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3721 = in0;
    end

    reg [7:0] out3722;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3722 = in0;
    end

    reg [7:0] out3723;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3723 = in0;
    end

    reg [7:0] out3724;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3724 = in0;
    end

    reg [7:0] out3725;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3725 = in0;
    end

    reg [7:0] out3726;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3726 = in0;
    end

    reg [7:0] out3727;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3727 = in0;
    end

    reg [7:0] out3728;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3728 = in0;
    end

    reg [7:0] out3729;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3729 = in0;
    end

    reg [7:0] out3730;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3730 = in0;
    end

    reg [7:0] out3731;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3731 = in0;
    end

    reg [7:0] out3732;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3732 = in0;
    end

    reg [7:0] out3733;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3733 = in0;
    end

    reg [7:0] out3734;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3734 = in0;
    end

    reg [7:0] out3735;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3735 = in0;
    end

    reg [7:0] out3736;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3736 = in0;
    end

    reg [7:0] out3737;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3737 = in0;
    end

    reg [7:0] out3738;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3738 = in0;
    end

    reg [7:0] out3739;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3739 = in0;
    end

    reg [7:0] out3740;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3740 = in0;
    end

    reg [7:0] out3741;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3741 = in0;
    end

    reg [7:0] out3742;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3742 = in0;
    end

    reg [7:0] out3743;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3743 = in0;
    end

    reg [7:0] out3744;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3744 = in0;
    end

    reg [7:0] out3745;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3745 = in0;
    end

    reg [7:0] out3746;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3746 = in0;
    end

    reg [7:0] out3747;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3747 = in0;
    end

    reg [7:0] out3748;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3748 = in0;
    end

    reg [7:0] out3749;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3749 = in0;
    end

    reg [7:0] out3750;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3750 = in0;
    end

    reg [7:0] out3751;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3751 = in0;
    end

    reg [7:0] out3752;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3752 = in0;
    end

    reg [7:0] out3753;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3753 = in0;
    end

    reg [7:0] out3754;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3754 = in0;
    end

    reg [7:0] out3755;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3755 = in0;
    end

    reg [7:0] out3756;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3756 = in0;
    end

    reg [7:0] out3757;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3757 = in0;
    end

    reg [7:0] out3758;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3758 = in0;
    end

    reg [7:0] out3759;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3759 = in0;
    end

    reg [7:0] out3760;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3760 = in0;
    end

    reg [7:0] out3761;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3761 = in0;
    end

    reg [7:0] out3762;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3762 = in0;
    end

    reg [7:0] out3763;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3763 = in0;
    end

    reg [7:0] out3764;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3764 = in0;
    end

    reg [7:0] out3765;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3765 = in0;
    end

    reg [7:0] out3766;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3766 = in0;
    end

    reg [7:0] out3767;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3767 = in0;
    end

    reg [7:0] out3768;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3768 = in0;
    end

    reg [7:0] out3769;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3769 = in0;
    end

    reg [7:0] out3770;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3770 = in0;
    end

    reg [7:0] out3771;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3771 = in0;
    end

    reg [7:0] out3772;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3772 = in0;
    end

    reg [7:0] out3773;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3773 = in0;
    end

    reg [7:0] out3774;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3774 = in0;
    end

    reg [7:0] out3775;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3775 = in0;
    end

    reg [7:0] out3776;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3776 = in0;
    end

    reg [7:0] out3777;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3777 = in0;
    end

    reg [7:0] out3778;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3778 = in0;
    end

    reg [7:0] out3779;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3779 = in0;
    end

    reg [7:0] out3780;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3780 = in0;
    end

    reg [7:0] out3781;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3781 = in0;
    end

    reg [7:0] out3782;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3782 = in0;
    end

    reg [7:0] out3783;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3783 = in0;
    end

    reg [7:0] out3784;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3784 = in0;
    end

    reg [7:0] out3785;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3785 = in0;
    end

    reg [7:0] out3786;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3786 = in0;
    end

    reg [7:0] out3787;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3787 = in0;
    end

    reg [7:0] out3788;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3788 = in0;
    end

    reg [7:0] out3789;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3789 = in0;
    end

    reg [7:0] out3790;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3790 = in0;
    end

    reg [7:0] out3791;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3791 = in0;
    end

    reg [7:0] out3792;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3792 = in0;
    end

    reg [7:0] out3793;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3793 = in0;
    end

    reg [7:0] out3794;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3794 = in0;
    end

    reg [7:0] out3795;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3795 = in0;
    end

    reg [7:0] out3796;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3796 = in0;
    end

    reg [7:0] out3797;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3797 = in0;
    end

    reg [7:0] out3798;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3798 = in0;
    end

    reg [7:0] out3799;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3799 = in0;
    end

    reg [7:0] out3800;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3800 = in0;
    end

    reg [7:0] out3801;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3801 = in0;
    end

    reg [7:0] out3802;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3802 = in0;
    end

    reg [7:0] out3803;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3803 = in0;
    end

    reg [7:0] out3804;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3804 = in0;
    end

    reg [7:0] out3805;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3805 = in0;
    end

    reg [7:0] out3806;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3806 = in0;
    end

    reg [7:0] out3807;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3807 = in0;
    end

    reg [7:0] out3808;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3808 = in0;
    end

    reg [7:0] out3809;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3809 = in0;
    end

    reg [7:0] out3810;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3810 = in0;
    end

    reg [7:0] out3811;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3811 = in0;
    end

    reg [7:0] out3812;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3812 = in0;
    end

    reg [7:0] out3813;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3813 = in0;
    end

    reg [7:0] out3814;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3814 = in0;
    end

    reg [7:0] out3815;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3815 = in0;
    end

    reg [7:0] out3816;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3816 = in0;
    end

    reg [7:0] out3817;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3817 = in0;
    end

    reg [7:0] out3818;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3818 = in0;
    end

    reg [7:0] out3819;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3819 = in0;
    end

    reg [7:0] out3820;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3820 = in0;
    end

    reg [7:0] out3821;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3821 = in0;
    end

    reg [7:0] out3822;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3822 = in0;
    end

    reg [7:0] out3823;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3823 = in0;
    end

    reg [7:0] out3824;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3824 = in0;
    end

    reg [7:0] out3825;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3825 = in0;
    end

    reg [7:0] out3826;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3826 = in0;
    end

    reg [7:0] out3827;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3827 = in0;
    end

    reg [7:0] out3828;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3828 = in0;
    end

    reg [7:0] out3829;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3829 = in0;
    end

    reg [7:0] out3830;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3830 = in0;
    end

    reg [7:0] out3831;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3831 = in0;
    end

    reg [7:0] out3832;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3832 = in0;
    end

    reg [7:0] out3833;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3833 = in0;
    end

    reg [7:0] out3834;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3834 = in0;
    end

    reg [7:0] out3835;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3835 = in0;
    end

    reg [7:0] out3836;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3836 = in0;
    end

    reg [7:0] out3837;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3837 = in0;
    end

    reg [7:0] out3838;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3838 = in0;
    end

    reg [7:0] out3839;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3839 = in0;
    end

    reg [7:0] out3840;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3840 = in0;
    end

    reg [7:0] out3841;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3841 = in0;
    end

    reg [7:0] out3842;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3842 = in0;
    end

    reg [7:0] out3843;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3843 = in0;
    end

    reg [7:0] out3844;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3844 = in0;
    end

    reg [7:0] out3845;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3845 = in0;
    end

    reg [7:0] out3846;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3846 = in0;
    end

    reg [7:0] out3847;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3847 = in0;
    end

    reg [7:0] out3848;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3848 = in0;
    end

    reg [7:0] out3849;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3849 = in0;
    end

    reg [7:0] out3850;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3850 = in0;
    end

    reg [7:0] out3851;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3851 = in0;
    end

    reg [7:0] out3852;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3852 = in0;
    end

    reg [7:0] out3853;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3853 = in0;
    end

    reg [7:0] out3854;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3854 = in0;
    end

    reg [7:0] out3855;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3855 = in0;
    end

    reg [7:0] out3856;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3856 = in0;
    end

    reg [7:0] out3857;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3857 = in0;
    end

    reg [7:0] out3858;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3858 = in0;
    end

    reg [7:0] out3859;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3859 = in0;
    end

    reg [7:0] out3860;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3860 = in0;
    end

    reg [7:0] out3861;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3861 = in0;
    end

    reg [7:0] out3862;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3862 = in0;
    end

    reg [7:0] out3863;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3863 = in0;
    end

    reg [7:0] out3864;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3864 = in0;
    end

    reg [7:0] out3865;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3865 = in0;
    end

    reg [7:0] out3866;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3866 = in0;
    end

    reg [7:0] out3867;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3867 = in0;
    end

    reg [7:0] out3868;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3868 = in0;
    end

    reg [7:0] out3869;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3869 = in0;
    end

    reg [7:0] out3870;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3870 = in0;
    end

    reg [7:0] out3871;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3871 = in0;
    end

    reg [7:0] out3872;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3872 = in0;
    end

    reg [7:0] out3873;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3873 = in0;
    end

    reg [7:0] out3874;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3874 = in0;
    end

    reg [7:0] out3875;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3875 = in0;
    end

    reg [7:0] out3876;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3876 = in0;
    end

    reg [7:0] out3877;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3877 = in0;
    end

    reg [7:0] out3878;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3878 = in0;
    end

    reg [7:0] out3879;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3879 = in0;
    end

    reg [7:0] out3880;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3880 = in0;
    end

    reg [7:0] out3881;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3881 = in0;
    end

    reg [7:0] out3882;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3882 = in0;
    end

    reg [7:0] out3883;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3883 = in0;
    end

    reg [7:0] out3884;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3884 = in0;
    end

    reg [7:0] out3885;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3885 = in0;
    end

    reg [7:0] out3886;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3886 = in0;
    end

    reg [7:0] out3887;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3887 = in0;
    end

    reg [7:0] out3888;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3888 = in0;
    end

    reg [7:0] out3889;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3889 = in0;
    end

    reg [7:0] out3890;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3890 = in0;
    end

    reg [7:0] out3891;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3891 = in0;
    end

    reg [7:0] out3892;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3892 = in0;
    end

    reg [7:0] out3893;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3893 = in0;
    end

    reg [7:0] out3894;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3894 = in0;
    end

    reg [7:0] out3895;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3895 = in0;
    end

    reg [7:0] out3896;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3896 = in0;
    end

    reg [7:0] out3897;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3897 = in0;
    end

    reg [7:0] out3898;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3898 = in0;
    end

    reg [7:0] out3899;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3899 = in0;
    end

    reg [7:0] out3900;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3900 = in0;
    end

    reg [7:0] out3901;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3901 = in0;
    end

    reg [7:0] out3902;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3902 = in0;
    end

    reg [7:0] out3903;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3903 = in0;
    end

    reg [7:0] out3904;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3904 = in0;
    end

    reg [7:0] out3905;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3905 = in0;
    end

    reg [7:0] out3906;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3906 = in0;
    end

    reg [7:0] out3907;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3907 = in0;
    end

    reg [7:0] out3908;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3908 = in0;
    end

    reg [7:0] out3909;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3909 = in0;
    end

    reg [7:0] out3910;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3910 = in0;
    end

    reg [7:0] out3911;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3911 = in0;
    end

    reg [7:0] out3912;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3912 = in0;
    end

    reg [7:0] out3913;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3913 = in0;
    end

    reg [7:0] out3914;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3914 = in0;
    end

    reg [7:0] out3915;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3915 = in0;
    end

    reg [7:0] out3916;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3916 = in0;
    end

    reg [7:0] out3917;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3917 = in0;
    end

    reg [7:0] out3918;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3918 = in0;
    end

    reg [7:0] out3919;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3919 = in0;
    end

    reg [7:0] out3920;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3920 = in0;
    end

    reg [7:0] out3921;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3921 = in0;
    end

    reg [7:0] out3922;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3922 = in0;
    end

    reg [7:0] out3923;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3923 = in0;
    end

    reg [7:0] out3924;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3924 = in0;
    end

    reg [7:0] out3925;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3925 = in0;
    end

    reg [7:0] out3926;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3926 = in0;
    end

    reg [7:0] out3927;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3927 = in0;
    end

    reg [7:0] out3928;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3928 = in0;
    end

    reg [7:0] out3929;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3929 = in0;
    end

    reg [7:0] out3930;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3930 = in0;
    end

    reg [7:0] out3931;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3931 = in0;
    end

    reg [7:0] out3932;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3932 = in0;
    end

    reg [7:0] out3933;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3933 = in0;
    end

    reg [7:0] out3934;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3934 = in0;
    end

    reg [7:0] out3935;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3935 = in0;
    end

    reg [7:0] out3936;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3936 = in0;
    end

    reg [7:0] out3937;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3937 = in0;
    end

    reg [7:0] out3938;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3938 = in0;
    end

    reg [7:0] out3939;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3939 = in0;
    end

    reg [7:0] out3940;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3940 = in0;
    end

    reg [7:0] out3941;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3941 = in0;
    end

    reg [7:0] out3942;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3942 = in0;
    end

    reg [7:0] out3943;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3943 = in0;
    end

    reg [7:0] out3944;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3944 = in0;
    end

    reg [7:0] out3945;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3945 = in0;
    end

    reg [7:0] out3946;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3946 = in0;
    end

    reg [7:0] out3947;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3947 = in0;
    end

    reg [7:0] out3948;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3948 = in0;
    end

    reg [7:0] out3949;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3949 = in0;
    end

    reg [7:0] out3950;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3950 = in0;
    end

    reg [7:0] out3951;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3951 = in0;
    end

    reg [7:0] out3952;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3952 = in0;
    end

    reg [7:0] out3953;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3953 = in0;
    end

    reg [7:0] out3954;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3954 = in0;
    end

    reg [7:0] out3955;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3955 = in0;
    end

    reg [7:0] out3956;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3956 = in0;
    end

    reg [7:0] out3957;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3957 = in0;
    end

    reg [7:0] out3958;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3958 = in0;
    end

    reg [7:0] out3959;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3959 = in0;
    end

    reg [7:0] out3960;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3960 = in0;
    end

    reg [7:0] out3961;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3961 = in0;
    end

    reg [7:0] out3962;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3962 = in0;
    end

    reg [7:0] out3963;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3963 = in0;
    end

    reg [7:0] out3964;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3964 = in0;
    end

    reg [7:0] out3965;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3965 = in0;
    end

    reg [7:0] out3966;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3966 = in0;
    end

    reg [7:0] out3967;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3967 = in0;
    end

    reg [7:0] out3968;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3968 = in0;
    end

    reg [7:0] out3969;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3969 = in0;
    end

    reg [7:0] out3970;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3970 = in0;
    end

    reg [7:0] out3971;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3971 = in0;
    end

    reg [7:0] out3972;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3972 = in0;
    end

    reg [7:0] out3973;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3973 = in0;
    end

    reg [7:0] out3974;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3974 = in0;
    end

    reg [7:0] out3975;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3975 = in0;
    end

    reg [7:0] out3976;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3976 = in0;
    end

    reg [7:0] out3977;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3977 = in0;
    end

    reg [7:0] out3978;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3978 = in0;
    end

    reg [7:0] out3979;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3979 = in0;
    end

    reg [7:0] out3980;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3980 = in0;
    end

    reg [7:0] out3981;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3981 = in0;
    end

    reg [7:0] out3982;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3982 = in0;
    end

    reg [7:0] out3983;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3983 = in0;
    end

    reg [7:0] out3984;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3984 = in0;
    end

    reg [7:0] out3985;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3985 = in0;
    end

    reg [7:0] out3986;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3986 = in0;
    end

    reg [7:0] out3987;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3987 = in0;
    end

    reg [7:0] out3988;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3988 = in0;
    end

    reg [7:0] out3989;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3989 = in0;
    end

    reg [7:0] out3990;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3990 = in0;
    end

    reg [7:0] out3991;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3991 = in0;
    end

    reg [7:0] out3992;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3992 = in0;
    end

    reg [7:0] out3993;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3993 = in0;
    end

    reg [7:0] out3994;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3994 = in0;
    end

    reg [7:0] out3995;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3995 = in0;
    end

    reg [7:0] out3996;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3996 = in0;
    end

    reg [7:0] out3997;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3997 = in0;
    end

    reg [7:0] out3998;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3998 = in0;
    end

    reg [7:0] out3999;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out3999 = in0;
    end

    reg [7:0] out4000;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4000 = in0;
    end

    reg [7:0] out4001;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4001 = in0;
    end

    reg [7:0] out4002;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4002 = in0;
    end

    reg [7:0] out4003;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4003 = in0;
    end

    reg [7:0] out4004;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4004 = in0;
    end

    reg [7:0] out4005;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4005 = in0;
    end

    reg [7:0] out4006;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4006 = in0;
    end

    reg [7:0] out4007;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4007 = in0;
    end

    reg [7:0] out4008;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4008 = in0;
    end

    reg [7:0] out4009;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4009 = in0;
    end

    reg [7:0] out4010;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4010 = in0;
    end

    reg [7:0] out4011;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4011 = in0;
    end

    reg [7:0] out4012;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4012 = in0;
    end

    reg [7:0] out4013;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4013 = in0;
    end

    reg [7:0] out4014;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4014 = in0;
    end

    reg [7:0] out4015;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4015 = in0;
    end

    reg [7:0] out4016;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4016 = in0;
    end

    reg [7:0] out4017;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4017 = in0;
    end

    reg [7:0] out4018;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4018 = in0;
    end

    reg [7:0] out4019;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4019 = in0;
    end

    reg [7:0] out4020;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4020 = in0;
    end

    reg [7:0] out4021;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4021 = in0;
    end

    reg [7:0] out4022;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4022 = in0;
    end

    reg [7:0] out4023;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4023 = in0;
    end

    reg [7:0] out4024;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4024 = in0;
    end

    reg [7:0] out4025;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4025 = in0;
    end

    reg [7:0] out4026;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4026 = in0;
    end

    reg [7:0] out4027;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4027 = in0;
    end

    reg [7:0] out4028;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4028 = in0;
    end

    reg [7:0] out4029;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4029 = in0;
    end

    reg [7:0] out4030;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4030 = in0;
    end

    reg [7:0] out4031;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4031 = in0;
    end

    reg [7:0] out4032;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4032 = in0;
    end

    reg [7:0] out4033;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4033 = in0;
    end

    reg [7:0] out4034;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4034 = in0;
    end

    reg [7:0] out4035;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4035 = in0;
    end

    reg [7:0] out4036;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4036 = in0;
    end

    reg [7:0] out4037;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4037 = in0;
    end

    reg [7:0] out4038;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4038 = in0;
    end

    reg [7:0] out4039;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4039 = in0;
    end

    reg [7:0] out4040;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4040 = in0;
    end

    reg [7:0] out4041;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4041 = in0;
    end

    reg [7:0] out4042;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4042 = in0;
    end

    reg [7:0] out4043;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4043 = in0;
    end

    reg [7:0] out4044;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4044 = in0;
    end

    reg [7:0] out4045;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4045 = in0;
    end

    reg [7:0] out4046;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4046 = in0;
    end

    reg [7:0] out4047;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4047 = in0;
    end

    reg [7:0] out4048;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4048 = in0;
    end

    reg [7:0] out4049;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4049 = in0;
    end

    reg [7:0] out4050;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4050 = in0;
    end

    reg [7:0] out4051;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4051 = in0;
    end

    reg [7:0] out4052;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4052 = in0;
    end

    reg [7:0] out4053;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4053 = in0;
    end

    reg [7:0] out4054;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4054 = in0;
    end

    reg [7:0] out4055;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4055 = in0;
    end

    reg [7:0] out4056;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4056 = in0;
    end

    reg [7:0] out4057;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4057 = in0;
    end

    reg [7:0] out4058;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4058 = in0;
    end

    reg [7:0] out4059;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4059 = in0;
    end

    reg [7:0] out4060;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4060 = in0;
    end

    reg [7:0] out4061;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4061 = in0;
    end

    reg [7:0] out4062;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4062 = in0;
    end

    reg [7:0] out4063;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4063 = in0;
    end

    reg [7:0] out4064;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4064 = in0;
    end

    reg [7:0] out4065;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4065 = in0;
    end

    reg [7:0] out4066;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4066 = in0;
    end

    reg [7:0] out4067;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4067 = in0;
    end

    reg [7:0] out4068;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4068 = in0;
    end

    reg [7:0] out4069;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4069 = in0;
    end

    reg [7:0] out4070;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4070 = in0;
    end

    reg [7:0] out4071;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4071 = in0;
    end

    reg [7:0] out4072;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4072 = in0;
    end

    reg [7:0] out4073;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4073 = in0;
    end

    reg [7:0] out4074;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4074 = in0;
    end

    reg [7:0] out4075;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4075 = in0;
    end

    reg [7:0] out4076;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4076 = in0;
    end

    reg [7:0] out4077;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4077 = in0;
    end

    reg [7:0] out4078;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4078 = in0;
    end

    reg [7:0] out4079;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4079 = in0;
    end

    reg [7:0] out4080;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4080 = in0;
    end

    reg [7:0] out4081;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4081 = in0;
    end

    reg [7:0] out4082;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4082 = in0;
    end

    reg [7:0] out4083;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4083 = in0;
    end

    reg [7:0] out4084;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4084 = in0;
    end

    reg [7:0] out4085;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4085 = in0;
    end

    reg [7:0] out4086;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4086 = in0;
    end

    reg [7:0] out4087;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4087 = in0;
    end

    reg [7:0] out4088;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4088 = in0;
    end

    reg [7:0] out4089;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4089 = in0;
    end

    reg [7:0] out4090;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4090 = in0;
    end

    reg [7:0] out4091;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4091 = in0;
    end

    reg [7:0] out4092;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4092 = in0;
    end

    reg [7:0] out4093;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4093 = in0;
    end

    reg [7:0] out4094;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4094 = in0;
    end

    reg [7:0] out4095;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4095 = in0;
    end

    reg [7:0] out4096;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4096 = in0;
    end

    reg [7:0] out4097;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4097 = in0;
    end

    reg [7:0] out4098;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4098 = in0;
    end

    reg [7:0] out4099;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4099 = in0;
    end

    reg [7:0] out4100;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4100 = in0;
    end

    reg [7:0] out4101;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4101 = in0;
    end

    reg [7:0] out4102;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4102 = in0;
    end

    reg [7:0] out4103;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4103 = in0;
    end

    reg [7:0] out4104;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4104 = in0;
    end

    reg [7:0] out4105;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4105 = in0;
    end

    reg [7:0] out4106;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4106 = in0;
    end

    reg [7:0] out4107;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4107 = in0;
    end

    reg [7:0] out4108;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4108 = in0;
    end

    reg [7:0] out4109;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4109 = in0;
    end

    reg [7:0] out4110;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4110 = in0;
    end

    reg [7:0] out4111;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4111 = in0;
    end

    reg [7:0] out4112;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4112 = in0;
    end

    reg [7:0] out4113;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4113 = in0;
    end

    reg [7:0] out4114;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4114 = in0;
    end

    reg [7:0] out4115;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4115 = in0;
    end

    reg [7:0] out4116;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4116 = in0;
    end

    reg [7:0] out4117;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4117 = in0;
    end

    reg [7:0] out4118;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4118 = in0;
    end

    reg [7:0] out4119;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4119 = in0;
    end

    reg [7:0] out4120;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4120 = in0;
    end

    reg [7:0] out4121;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4121 = in0;
    end

    reg [7:0] out4122;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4122 = in0;
    end

    reg [7:0] out4123;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4123 = in0;
    end

    reg [7:0] out4124;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4124 = in0;
    end

    reg [7:0] out4125;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4125 = in0;
    end

    reg [7:0] out4126;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4126 = in0;
    end

    reg [7:0] out4127;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4127 = in0;
    end

    reg [7:0] out4128;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4128 = in0;
    end

    reg [7:0] out4129;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4129 = in0;
    end

    reg [7:0] out4130;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4130 = in0;
    end

    reg [7:0] out4131;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4131 = in0;
    end

    reg [7:0] out4132;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4132 = in0;
    end

    reg [7:0] out4133;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4133 = in0;
    end

    reg [7:0] out4134;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4134 = in0;
    end

    reg [7:0] out4135;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4135 = in0;
    end

    reg [7:0] out4136;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4136 = in0;
    end

    reg [7:0] out4137;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4137 = in0;
    end

    reg [7:0] out4138;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4138 = in0;
    end

    reg [7:0] out4139;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4139 = in0;
    end

    reg [7:0] out4140;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4140 = in0;
    end

    reg [7:0] out4141;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4141 = in0;
    end

    reg [7:0] out4142;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4142 = in0;
    end

    reg [7:0] out4143;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4143 = in0;
    end

    reg [7:0] out4144;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4144 = in0;
    end

    reg [7:0] out4145;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4145 = in0;
    end

    reg [7:0] out4146;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4146 = in0;
    end

    reg [7:0] out4147;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4147 = in0;
    end

    reg [7:0] out4148;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4148 = in0;
    end

    reg [7:0] out4149;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4149 = in0;
    end

    reg [7:0] out4150;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4150 = in0;
    end

    reg [7:0] out4151;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4151 = in0;
    end

    reg [7:0] out4152;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4152 = in0;
    end

    reg [7:0] out4153;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4153 = in0;
    end

    reg [7:0] out4154;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4154 = in0;
    end

    reg [7:0] out4155;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4155 = in0;
    end

    reg [7:0] out4156;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4156 = in0;
    end

    reg [7:0] out4157;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4157 = in0;
    end

    reg [7:0] out4158;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4158 = in0;
    end

    reg [7:0] out4159;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4159 = in0;
    end

    reg [7:0] out4160;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4160 = in0;
    end

    reg [7:0] out4161;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4161 = in0;
    end

    reg [7:0] out4162;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4162 = in0;
    end

    reg [7:0] out4163;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4163 = in0;
    end

    reg [7:0] out4164;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4164 = in0;
    end

    reg [7:0] out4165;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4165 = in0;
    end

    reg [7:0] out4166;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4166 = in0;
    end

    reg [7:0] out4167;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4167 = in0;
    end

    reg [7:0] out4168;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4168 = in0;
    end

    reg [7:0] out4169;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4169 = in0;
    end

    reg [7:0] out4170;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4170 = in0;
    end

    reg [7:0] out4171;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4171 = in0;
    end

    reg [7:0] out4172;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4172 = in0;
    end

    reg [7:0] out4173;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4173 = in0;
    end

    reg [7:0] out4174;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4174 = in0;
    end

    reg [7:0] out4175;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4175 = in0;
    end

    reg [7:0] out4176;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4176 = in0;
    end

    reg [7:0] out4177;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4177 = in0;
    end

    reg [7:0] out4178;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4178 = in0;
    end

    reg [7:0] out4179;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4179 = in0;
    end

    reg [7:0] out4180;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4180 = in0;
    end

    reg [7:0] out4181;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4181 = in0;
    end

    reg [7:0] out4182;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4182 = in0;
    end

    reg [7:0] out4183;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4183 = in0;
    end

    reg [7:0] out4184;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4184 = in0;
    end

    reg [7:0] out4185;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4185 = in0;
    end

    reg [7:0] out4186;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4186 = in0;
    end

    reg [7:0] out4187;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4187 = in0;
    end

    reg [7:0] out4188;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4188 = in0;
    end

    reg [7:0] out4189;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4189 = in0;
    end

    reg [7:0] out4190;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4190 = in0;
    end

    reg [7:0] out4191;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4191 = in0;
    end

    reg [7:0] out4192;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4192 = in0;
    end

    reg [7:0] out4193;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4193 = in0;
    end

    reg [7:0] out4194;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4194 = in0;
    end

    reg [7:0] out4195;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4195 = in0;
    end

    reg [7:0] out4196;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4196 = in0;
    end

    reg [7:0] out4197;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4197 = in0;
    end

    reg [7:0] out4198;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4198 = in0;
    end

    reg [7:0] out4199;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4199 = in0;
    end

    reg [7:0] out4200;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4200 = in0;
    end

    reg [7:0] out4201;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4201 = in0;
    end

    reg [7:0] out4202;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4202 = in0;
    end

    reg [7:0] out4203;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4203 = in0;
    end

    reg [7:0] out4204;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4204 = in0;
    end

    reg [7:0] out4205;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4205 = in0;
    end

    reg [7:0] out4206;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4206 = in0;
    end

    reg [7:0] out4207;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4207 = in0;
    end

    reg [7:0] out4208;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4208 = in0;
    end

    reg [7:0] out4209;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4209 = in0;
    end

    reg [7:0] out4210;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4210 = in0;
    end

    reg [7:0] out4211;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4211 = in0;
    end

    reg [7:0] out4212;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4212 = in0;
    end

    reg [7:0] out4213;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4213 = in0;
    end

    reg [7:0] out4214;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4214 = in0;
    end

    reg [7:0] out4215;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4215 = in0;
    end

    reg [7:0] out4216;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4216 = in0;
    end

    reg [7:0] out4217;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4217 = in0;
    end

    reg [7:0] out4218;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4218 = in0;
    end

    reg [7:0] out4219;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4219 = in0;
    end

    reg [7:0] out4220;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4220 = in0;
    end

    reg [7:0] out4221;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4221 = in0;
    end

    reg [7:0] out4222;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4222 = in0;
    end

    reg [7:0] out4223;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4223 = in0;
    end

    reg [7:0] out4224;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4224 = in0;
    end

    reg [7:0] out4225;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4225 = in0;
    end

    reg [7:0] out4226;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4226 = in0;
    end

    reg [7:0] out4227;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4227 = in0;
    end

    reg [7:0] out4228;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4228 = in0;
    end

    reg [7:0] out4229;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4229 = in0;
    end

    reg [7:0] out4230;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4230 = in0;
    end

    reg [7:0] out4231;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4231 = in0;
    end

    reg [7:0] out4232;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4232 = in0;
    end

    reg [7:0] out4233;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4233 = in0;
    end

    reg [7:0] out4234;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4234 = in0;
    end

    reg [7:0] out4235;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4235 = in0;
    end

    reg [7:0] out4236;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4236 = in0;
    end

    reg [7:0] out4237;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4237 = in0;
    end

    reg [7:0] out4238;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4238 = in0;
    end

    reg [7:0] out4239;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4239 = in0;
    end

    reg [7:0] out4240;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4240 = in0;
    end

    reg [7:0] out4241;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4241 = in0;
    end

    reg [7:0] out4242;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4242 = in0;
    end

    reg [7:0] out4243;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4243 = in0;
    end

    reg [7:0] out4244;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4244 = in0;
    end

    reg [7:0] out4245;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4245 = in0;
    end

    reg [7:0] out4246;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4246 = in0;
    end

    reg [7:0] out4247;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4247 = in0;
    end

    reg [7:0] out4248;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4248 = in0;
    end

    reg [7:0] out4249;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4249 = in0;
    end

    reg [7:0] out4250;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4250 = in0;
    end

    reg [7:0] out4251;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4251 = in0;
    end

    reg [7:0] out4252;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4252 = in0;
    end

    reg [7:0] out4253;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4253 = in0;
    end

    reg [7:0] out4254;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4254 = in0;
    end

    reg [7:0] out4255;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4255 = in0;
    end

    reg [7:0] out4256;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4256 = in0;
    end

    reg [7:0] out4257;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4257 = in0;
    end

    reg [7:0] out4258;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4258 = in0;
    end

    reg [7:0] out4259;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4259 = in0;
    end

    reg [7:0] out4260;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4260 = in0;
    end

    reg [7:0] out4261;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4261 = in0;
    end

    reg [7:0] out4262;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4262 = in0;
    end

    reg [7:0] out4263;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4263 = in0;
    end

    reg [7:0] out4264;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4264 = in0;
    end

    reg [7:0] out4265;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4265 = in0;
    end

    reg [7:0] out4266;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4266 = in0;
    end

    reg [7:0] out4267;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4267 = in0;
    end

    reg [7:0] out4268;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4268 = in0;
    end

    reg [7:0] out4269;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4269 = in0;
    end

    reg [7:0] out4270;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4270 = in0;
    end

    reg [7:0] out4271;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4271 = in0;
    end

    reg [7:0] out4272;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4272 = in0;
    end

    reg [7:0] out4273;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4273 = in0;
    end

    reg [7:0] out4274;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4274 = in0;
    end

    reg [7:0] out4275;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4275 = in0;
    end

    reg [7:0] out4276;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4276 = in0;
    end

    reg [7:0] out4277;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4277 = in0;
    end

    reg [7:0] out4278;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4278 = in0;
    end

    reg [7:0] out4279;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4279 = in0;
    end

    reg [7:0] out4280;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4280 = in0;
    end

    reg [7:0] out4281;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4281 = in0;
    end

    reg [7:0] out4282;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4282 = in0;
    end

    reg [7:0] out4283;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4283 = in0;
    end

    reg [7:0] out4284;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4284 = in0;
    end

    reg [7:0] out4285;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4285 = in0;
    end

    reg [7:0] out4286;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4286 = in0;
    end

    reg [7:0] out4287;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4287 = in0;
    end

    reg [7:0] out4288;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4288 = in0;
    end

    reg [7:0] out4289;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4289 = in0;
    end

    reg [7:0] out4290;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4290 = in0;
    end

    reg [7:0] out4291;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4291 = in0;
    end

    reg [7:0] out4292;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4292 = in0;
    end

    reg [7:0] out4293;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4293 = in0;
    end

    reg [7:0] out4294;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4294 = in0;
    end

    reg [7:0] out4295;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4295 = in0;
    end

    reg [7:0] out4296;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4296 = in0;
    end

    reg [7:0] out4297;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4297 = in0;
    end

    reg [7:0] out4298;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4298 = in0;
    end

    reg [7:0] out4299;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4299 = in0;
    end

    reg [7:0] out4300;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4300 = in0;
    end

    reg [7:0] out4301;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4301 = in0;
    end

    reg [7:0] out4302;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4302 = in0;
    end

    reg [7:0] out4303;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4303 = in0;
    end

    reg [7:0] out4304;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4304 = in0;
    end

    reg [7:0] out4305;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4305 = in0;
    end

    reg [7:0] out4306;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4306 = in0;
    end

    reg [7:0] out4307;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4307 = in0;
    end

    reg [7:0] out4308;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4308 = in0;
    end

    reg [7:0] out4309;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4309 = in0;
    end

    reg [7:0] out4310;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4310 = in0;
    end

    reg [7:0] out4311;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4311 = in0;
    end

    reg [7:0] out4312;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4312 = in0;
    end

    reg [7:0] out4313;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4313 = in0;
    end

    reg [7:0] out4314;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4314 = in0;
    end

    reg [7:0] out4315;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4315 = in0;
    end

    reg [7:0] out4316;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4316 = in0;
    end

    reg [7:0] out4317;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4317 = in0;
    end

    reg [7:0] out4318;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4318 = in0;
    end

    reg [7:0] out4319;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4319 = in0;
    end

    reg [7:0] out4320;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4320 = in0;
    end

    reg [7:0] out4321;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4321 = in0;
    end

    reg [7:0] out4322;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4322 = in0;
    end

    reg [7:0] out4323;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4323 = in0;
    end

    reg [7:0] out4324;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4324 = in0;
    end

    reg [7:0] out4325;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4325 = in0;
    end

    reg [7:0] out4326;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4326 = in0;
    end

    reg [7:0] out4327;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4327 = in0;
    end

    reg [7:0] out4328;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4328 = in0;
    end

    reg [7:0] out4329;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4329 = in0;
    end

    reg [7:0] out4330;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4330 = in0;
    end

    reg [7:0] out4331;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4331 = in0;
    end

    reg [7:0] out4332;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4332 = in0;
    end

    reg [7:0] out4333;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4333 = in0;
    end

    reg [7:0] out4334;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4334 = in0;
    end

    reg [7:0] out4335;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4335 = in0;
    end

    reg [7:0] out4336;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4336 = in0;
    end

    reg [7:0] out4337;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4337 = in0;
    end

    reg [7:0] out4338;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4338 = in0;
    end

    reg [7:0] out4339;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4339 = in0;
    end

    reg [7:0] out4340;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4340 = in0;
    end

    reg [7:0] out4341;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4341 = in0;
    end

    reg [7:0] out4342;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4342 = in0;
    end

    reg [7:0] out4343;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4343 = in0;
    end

    reg [7:0] out4344;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4344 = in0;
    end

    reg [7:0] out4345;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4345 = in0;
    end

    reg [7:0] out4346;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4346 = in0;
    end

    reg [7:0] out4347;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4347 = in0;
    end

    reg [7:0] out4348;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4348 = in0;
    end

    reg [7:0] out4349;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4349 = in0;
    end

    reg [7:0] out4350;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4350 = in0;
    end

    reg [7:0] out4351;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4351 = in0;
    end

    reg [7:0] out4352;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4352 = in0;
    end

    reg [7:0] out4353;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4353 = in0;
    end

    reg [7:0] out4354;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4354 = in0;
    end

    reg [7:0] out4355;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4355 = in0;
    end

    reg [7:0] out4356;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4356 = in0;
    end

    reg [7:0] out4357;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4357 = in0;
    end

    reg [7:0] out4358;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4358 = in0;
    end

    reg [7:0] out4359;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4359 = in0;
    end

    reg [7:0] out4360;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4360 = in0;
    end

    reg [7:0] out4361;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4361 = in0;
    end

    reg [7:0] out4362;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4362 = in0;
    end

    reg [7:0] out4363;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4363 = in0;
    end

    reg [7:0] out4364;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4364 = in0;
    end

    reg [7:0] out4365;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4365 = in0;
    end

    reg [7:0] out4366;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4366 = in0;
    end

    reg [7:0] out4367;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4367 = in0;
    end

    reg [7:0] out4368;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4368 = in0;
    end

    reg [7:0] out4369;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4369 = in0;
    end

    reg [7:0] out4370;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4370 = in0;
    end

    reg [7:0] out4371;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4371 = in0;
    end

    reg [7:0] out4372;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4372 = in0;
    end

    reg [7:0] out4373;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4373 = in0;
    end

    reg [7:0] out4374;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4374 = in0;
    end

    reg [7:0] out4375;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4375 = in0;
    end

    reg [7:0] out4376;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4376 = in0;
    end

    reg [7:0] out4377;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4377 = in0;
    end

    reg [7:0] out4378;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4378 = in0;
    end

    reg [7:0] out4379;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4379 = in0;
    end

    reg [7:0] out4380;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4380 = in0;
    end

    reg [7:0] out4381;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4381 = in0;
    end

    reg [7:0] out4382;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4382 = in0;
    end

    reg [7:0] out4383;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4383 = in0;
    end

    reg [7:0] out4384;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4384 = in0;
    end

    reg [7:0] out4385;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4385 = in0;
    end

    reg [7:0] out4386;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4386 = in0;
    end

    reg [7:0] out4387;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4387 = in0;
    end

    reg [7:0] out4388;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4388 = in0;
    end

    reg [7:0] out4389;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4389 = in0;
    end

    reg [7:0] out4390;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4390 = in0;
    end

    reg [7:0] out4391;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4391 = in0;
    end

    reg [7:0] out4392;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4392 = in0;
    end

    reg [7:0] out4393;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4393 = in0;
    end

    reg [7:0] out4394;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4394 = in0;
    end

    reg [7:0] out4395;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4395 = in0;
    end

    reg [7:0] out4396;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4396 = in0;
    end

    reg [7:0] out4397;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4397 = in0;
    end

    reg [7:0] out4398;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4398 = in0;
    end

    reg [7:0] out4399;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4399 = in0;
    end

    reg [7:0] out4400;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4400 = in0;
    end

    reg [7:0] out4401;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4401 = in0;
    end

    reg [7:0] out4402;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4402 = in0;
    end

    reg [7:0] out4403;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4403 = in0;
    end

    reg [7:0] out4404;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4404 = in0;
    end

    reg [7:0] out4405;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4405 = in0;
    end

    reg [7:0] out4406;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4406 = in0;
    end

    reg [7:0] out4407;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4407 = in0;
    end

    reg [7:0] out4408;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4408 = in0;
    end

    reg [7:0] out4409;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4409 = in0;
    end

    reg [7:0] out4410;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4410 = in0;
    end

    reg [7:0] out4411;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4411 = in0;
    end

    reg [7:0] out4412;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4412 = in0;
    end

    reg [7:0] out4413;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4413 = in0;
    end

    reg [7:0] out4414;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4414 = in0;
    end

    reg [7:0] out4415;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4415 = in0;
    end

    reg [7:0] out4416;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4416 = in0;
    end

    reg [7:0] out4417;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4417 = in0;
    end

    reg [7:0] out4418;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4418 = in0;
    end

    reg [7:0] out4419;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4419 = in0;
    end

    reg [7:0] out4420;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4420 = in0;
    end

    reg [7:0] out4421;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4421 = in0;
    end

    reg [7:0] out4422;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4422 = in0;
    end

    reg [7:0] out4423;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4423 = in0;
    end

    reg [7:0] out4424;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4424 = in0;
    end

    reg [7:0] out4425;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4425 = in0;
    end

    reg [7:0] out4426;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4426 = in0;
    end

    reg [7:0] out4427;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4427 = in0;
    end

    reg [7:0] out4428;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4428 = in0;
    end

    reg [7:0] out4429;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4429 = in0;
    end

    reg [7:0] out4430;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4430 = in0;
    end

    reg [7:0] out4431;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4431 = in0;
    end

    reg [7:0] out4432;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4432 = in0;
    end

    reg [7:0] out4433;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4433 = in0;
    end

    reg [7:0] out4434;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4434 = in0;
    end

    reg [7:0] out4435;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4435 = in0;
    end

    reg [7:0] out4436;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4436 = in0;
    end

    reg [7:0] out4437;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4437 = in0;
    end

    reg [7:0] out4438;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4438 = in0;
    end

    reg [7:0] out4439;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4439 = in0;
    end

    reg [7:0] out4440;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4440 = in0;
    end

    reg [7:0] out4441;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4441 = in0;
    end

    reg [7:0] out4442;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4442 = in0;
    end

    reg [7:0] out4443;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4443 = in0;
    end

    reg [7:0] out4444;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4444 = in0;
    end

    reg [7:0] out4445;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4445 = in0;
    end

    reg [7:0] out4446;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4446 = in0;
    end

    reg [7:0] out4447;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4447 = in0;
    end

    reg [7:0] out4448;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4448 = in0;
    end

    reg [7:0] out4449;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4449 = in0;
    end

    reg [7:0] out4450;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4450 = in0;
    end

    reg [7:0] out4451;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4451 = in0;
    end

    reg [7:0] out4452;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4452 = in0;
    end

    reg [7:0] out4453;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4453 = in0;
    end

    reg [7:0] out4454;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4454 = in0;
    end

    reg [7:0] out4455;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4455 = in0;
    end

    reg [7:0] out4456;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4456 = in0;
    end

    reg [7:0] out4457;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4457 = in0;
    end

    reg [7:0] out4458;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4458 = in0;
    end

    reg [7:0] out4459;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4459 = in0;
    end

    reg [7:0] out4460;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4460 = in0;
    end

    reg [7:0] out4461;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4461 = in0;
    end

    reg [7:0] out4462;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4462 = in0;
    end

    reg [7:0] out4463;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4463 = in0;
    end

    reg [7:0] out4464;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4464 = in0;
    end

    reg [7:0] out4465;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4465 = in0;
    end

    reg [7:0] out4466;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4466 = in0;
    end

    reg [7:0] out4467;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4467 = in0;
    end

    reg [7:0] out4468;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4468 = in0;
    end

    reg [7:0] out4469;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4469 = in0;
    end

    reg [7:0] out4470;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4470 = in0;
    end

    reg [7:0] out4471;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4471 = in0;
    end

    reg [7:0] out4472;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4472 = in0;
    end

    reg [7:0] out4473;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4473 = in0;
    end

    reg [7:0] out4474;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4474 = in0;
    end

    reg [7:0] out4475;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4475 = in0;
    end

    reg [7:0] out4476;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4476 = in0;
    end

    reg [7:0] out4477;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4477 = in0;
    end

    reg [7:0] out4478;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4478 = in0;
    end

    reg [7:0] out4479;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4479 = in0;
    end

    reg [7:0] out4480;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4480 = in0;
    end

    reg [7:0] out4481;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4481 = in0;
    end

    reg [7:0] out4482;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4482 = in0;
    end

    reg [7:0] out4483;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4483 = in0;
    end

    reg [7:0] out4484;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4484 = in0;
    end

    reg [7:0] out4485;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4485 = in0;
    end

    reg [7:0] out4486;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4486 = in0;
    end

    reg [7:0] out4487;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4487 = in0;
    end

    reg [7:0] out4488;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4488 = in0;
    end

    reg [7:0] out4489;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4489 = in0;
    end

    reg [7:0] out4490;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4490 = in0;
    end

    reg [7:0] out4491;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4491 = in0;
    end

    reg [7:0] out4492;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4492 = in0;
    end

    reg [7:0] out4493;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4493 = in0;
    end

    reg [7:0] out4494;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4494 = in0;
    end

    reg [7:0] out4495;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4495 = in0;
    end

    reg [7:0] out4496;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4496 = in0;
    end

    reg [7:0] out4497;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4497 = in0;
    end

    reg [7:0] out4498;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4498 = in0;
    end

    reg [7:0] out4499;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4499 = in0;
    end

    reg [7:0] out4500;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4500 = in0;
    end

    reg [7:0] out4501;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4501 = in0;
    end

    reg [7:0] out4502;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4502 = in0;
    end

    reg [7:0] out4503;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4503 = in0;
    end

    reg [7:0] out4504;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4504 = in0;
    end

    reg [7:0] out4505;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4505 = in0;
    end

    reg [7:0] out4506;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4506 = in0;
    end

    reg [7:0] out4507;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4507 = in0;
    end

    reg [7:0] out4508;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4508 = in0;
    end

    reg [7:0] out4509;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4509 = in0;
    end

    reg [7:0] out4510;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4510 = in0;
    end

    reg [7:0] out4511;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4511 = in0;
    end

    reg [7:0] out4512;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4512 = in0;
    end

    reg [7:0] out4513;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4513 = in0;
    end

    reg [7:0] out4514;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4514 = in0;
    end

    reg [7:0] out4515;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4515 = in0;
    end

    reg [7:0] out4516;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4516 = in0;
    end

    reg [7:0] out4517;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4517 = in0;
    end

    reg [7:0] out4518;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4518 = in0;
    end

    reg [7:0] out4519;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4519 = in0;
    end

    reg [7:0] out4520;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4520 = in0;
    end

    reg [7:0] out4521;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4521 = in0;
    end

    reg [7:0] out4522;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4522 = in0;
    end

    reg [7:0] out4523;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4523 = in0;
    end

    reg [7:0] out4524;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4524 = in0;
    end

    reg [7:0] out4525;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4525 = in0;
    end

    reg [7:0] out4526;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4526 = in0;
    end

    reg [7:0] out4527;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4527 = in0;
    end

    reg [7:0] out4528;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4528 = in0;
    end

    reg [7:0] out4529;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4529 = in0;
    end

    reg [7:0] out4530;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4530 = in0;
    end

    reg [7:0] out4531;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4531 = in0;
    end

    reg [7:0] out4532;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4532 = in0;
    end

    reg [7:0] out4533;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4533 = in0;
    end

    reg [7:0] out4534;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4534 = in0;
    end

    reg [7:0] out4535;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4535 = in0;
    end

    reg [7:0] out4536;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4536 = in0;
    end

    reg [7:0] out4537;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4537 = in0;
    end

    reg [7:0] out4538;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4538 = in0;
    end

    reg [7:0] out4539;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4539 = in0;
    end

    reg [7:0] out4540;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4540 = in0;
    end

    reg [7:0] out4541;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4541 = in0;
    end

    reg [7:0] out4542;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4542 = in0;
    end

    reg [7:0] out4543;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4543 = in0;
    end

    reg [7:0] out4544;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4544 = in0;
    end

    reg [7:0] out4545;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4545 = in0;
    end

    reg [7:0] out4546;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4546 = in0;
    end

    reg [7:0] out4547;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4547 = in0;
    end

    reg [7:0] out4548;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4548 = in0;
    end

    reg [7:0] out4549;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4549 = in0;
    end

    reg [7:0] out4550;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4550 = in0;
    end

    reg [7:0] out4551;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4551 = in0;
    end

    reg [7:0] out4552;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4552 = in0;
    end

    reg [7:0] out4553;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4553 = in0;
    end

    reg [7:0] out4554;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4554 = in0;
    end

    reg [7:0] out4555;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4555 = in0;
    end

    reg [7:0] out4556;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4556 = in0;
    end

    reg [7:0] out4557;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4557 = in0;
    end

    reg [7:0] out4558;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4558 = in0;
    end

    reg [7:0] out4559;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4559 = in0;
    end

    reg [7:0] out4560;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4560 = in0;
    end

    reg [7:0] out4561;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4561 = in0;
    end

    reg [7:0] out4562;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4562 = in0;
    end

    reg [7:0] out4563;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4563 = in0;
    end

    reg [7:0] out4564;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4564 = in0;
    end

    reg [7:0] out4565;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4565 = in0;
    end

    reg [7:0] out4566;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4566 = in0;
    end

    reg [7:0] out4567;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4567 = in0;
    end

    reg [7:0] out4568;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4568 = in0;
    end

    reg [7:0] out4569;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4569 = in0;
    end

    reg [7:0] out4570;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4570 = in0;
    end

    reg [7:0] out4571;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4571 = in0;
    end

    reg [7:0] out4572;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4572 = in0;
    end

    reg [7:0] out4573;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4573 = in0;
    end

    reg [7:0] out4574;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4574 = in0;
    end

    reg [7:0] out4575;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4575 = in0;
    end

    reg [7:0] out4576;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4576 = in0;
    end

    reg [7:0] out4577;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4577 = in0;
    end

    reg [7:0] out4578;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4578 = in0;
    end

    reg [7:0] out4579;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4579 = in0;
    end

    reg [7:0] out4580;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4580 = in0;
    end

    reg [7:0] out4581;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4581 = in0;
    end

    reg [7:0] out4582;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4582 = in0;
    end

    reg [7:0] out4583;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4583 = in0;
    end

    reg [7:0] out4584;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4584 = in0;
    end

    reg [7:0] out4585;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4585 = in0;
    end

    reg [7:0] out4586;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4586 = in0;
    end

    reg [7:0] out4587;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4587 = in0;
    end

    reg [7:0] out4588;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4588 = in0;
    end

    reg [7:0] out4589;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4589 = in0;
    end

    reg [7:0] out4590;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4590 = in0;
    end

    reg [7:0] out4591;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4591 = in0;
    end

    reg [7:0] out4592;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4592 = in0;
    end

    reg [7:0] out4593;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4593 = in0;
    end

    reg [7:0] out4594;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4594 = in0;
    end

    reg [7:0] out4595;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4595 = in0;
    end

    reg [7:0] out4596;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4596 = in0;
    end

    reg [7:0] out4597;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4597 = in0;
    end

    reg [7:0] out4598;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4598 = in0;
    end

    reg [7:0] out4599;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4599 = in0;
    end

    reg [7:0] out4600;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4600 = in0;
    end

    reg [7:0] out4601;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4601 = in0;
    end

    reg [7:0] out4602;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4602 = in0;
    end

    reg [7:0] out4603;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4603 = in0;
    end

    reg [7:0] out4604;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4604 = in0;
    end

    reg [7:0] out4605;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4605 = in0;
    end

    reg [7:0] out4606;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4606 = in0;
    end

    reg [7:0] out4607;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4607 = in0;
    end

    reg [7:0] out4608;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4608 = in0;
    end

    reg [7:0] out4609;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4609 = in0;
    end

    reg [7:0] out4610;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4610 = in0;
    end

    reg [7:0] out4611;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4611 = in0;
    end

    reg [7:0] out4612;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4612 = in0;
    end

    reg [7:0] out4613;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4613 = in0;
    end

    reg [7:0] out4614;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4614 = in0;
    end

    reg [7:0] out4615;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4615 = in0;
    end

    reg [7:0] out4616;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4616 = in0;
    end

    reg [7:0] out4617;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4617 = in0;
    end

    reg [7:0] out4618;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4618 = in0;
    end

    reg [7:0] out4619;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4619 = in0;
    end

    reg [7:0] out4620;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4620 = in0;
    end

    reg [7:0] out4621;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4621 = in0;
    end

    reg [7:0] out4622;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4622 = in0;
    end

    reg [7:0] out4623;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4623 = in0;
    end

    reg [7:0] out4624;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4624 = in0;
    end

    reg [7:0] out4625;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4625 = in0;
    end

    reg [7:0] out4626;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4626 = in0;
    end

    reg [7:0] out4627;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4627 = in0;
    end

    reg [7:0] out4628;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4628 = in0;
    end

    reg [7:0] out4629;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4629 = in0;
    end

    reg [7:0] out4630;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4630 = in0;
    end

    reg [7:0] out4631;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4631 = in0;
    end

    reg [7:0] out4632;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4632 = in0;
    end

    reg [7:0] out4633;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4633 = in0;
    end

    reg [7:0] out4634;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4634 = in0;
    end

    reg [7:0] out4635;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4635 = in0;
    end

    reg [7:0] out4636;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4636 = in0;
    end

    reg [7:0] out4637;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4637 = in0;
    end

    reg [7:0] out4638;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4638 = in0;
    end

    reg [7:0] out4639;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4639 = in0;
    end

    reg [7:0] out4640;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4640 = in0;
    end

    reg [7:0] out4641;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4641 = in0;
    end

    reg [7:0] out4642;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4642 = in0;
    end

    reg [7:0] out4643;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4643 = in0;
    end

    reg [7:0] out4644;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4644 = in0;
    end

    reg [7:0] out4645;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4645 = in0;
    end

    reg [7:0] out4646;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4646 = in0;
    end

    reg [7:0] out4647;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4647 = in0;
    end

    reg [7:0] out4648;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4648 = in0;
    end

    reg [7:0] out4649;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4649 = in0;
    end

    reg [7:0] out4650;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4650 = in0;
    end

    reg [7:0] out4651;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4651 = in0;
    end

    reg [7:0] out4652;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4652 = in0;
    end

    reg [7:0] out4653;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4653 = in0;
    end

    reg [7:0] out4654;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4654 = in0;
    end

    reg [7:0] out4655;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4655 = in0;
    end

    reg [7:0] out4656;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4656 = in0;
    end

    reg [7:0] out4657;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4657 = in0;
    end

    reg [7:0] out4658;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4658 = in0;
    end

    reg [7:0] out4659;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4659 = in0;
    end

    reg [7:0] out4660;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4660 = in0;
    end

    reg [7:0] out4661;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4661 = in0;
    end

    reg [7:0] out4662;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4662 = in0;
    end

    reg [7:0] out4663;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4663 = in0;
    end

    reg [7:0] out4664;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4664 = in0;
    end

    reg [7:0] out4665;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4665 = in0;
    end

    reg [7:0] out4666;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4666 = in0;
    end

    reg [7:0] out4667;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4667 = in0;
    end

    reg [7:0] out4668;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4668 = in0;
    end

    reg [7:0] out4669;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4669 = in0;
    end

    reg [7:0] out4670;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4670 = in0;
    end

    reg [7:0] out4671;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4671 = in0;
    end

    reg [7:0] out4672;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4672 = in0;
    end

    reg [7:0] out4673;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4673 = in0;
    end

    reg [7:0] out4674;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4674 = in0;
    end

    reg [7:0] out4675;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4675 = in0;
    end

    reg [7:0] out4676;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4676 = in0;
    end

    reg [7:0] out4677;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4677 = in0;
    end

    reg [7:0] out4678;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4678 = in0;
    end

    reg [7:0] out4679;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4679 = in0;
    end

    reg [7:0] out4680;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4680 = in0;
    end

    reg [7:0] out4681;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4681 = in0;
    end

    reg [7:0] out4682;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4682 = in0;
    end

    reg [7:0] out4683;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4683 = in0;
    end

    reg [7:0] out4684;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4684 = in0;
    end

    reg [7:0] out4685;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4685 = in0;
    end

    reg [7:0] out4686;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4686 = in0;
    end

    reg [7:0] out4687;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4687 = in0;
    end

    reg [7:0] out4688;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4688 = in0;
    end

    reg [7:0] out4689;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4689 = in0;
    end

    reg [7:0] out4690;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4690 = in0;
    end

    reg [7:0] out4691;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4691 = in0;
    end

    reg [7:0] out4692;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4692 = in0;
    end

    reg [7:0] out4693;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4693 = in0;
    end

    reg [7:0] out4694;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4694 = in0;
    end

    reg [7:0] out4695;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4695 = in0;
    end

    reg [7:0] out4696;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4696 = in0;
    end

    reg [7:0] out4697;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4697 = in0;
    end

    reg [7:0] out4698;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4698 = in0;
    end

    reg [7:0] out4699;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4699 = in0;
    end

    reg [7:0] out4700;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4700 = in0;
    end

    reg [7:0] out4701;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4701 = in0;
    end

    reg [7:0] out4702;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4702 = in0;
    end

    reg [7:0] out4703;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4703 = in0;
    end

    reg [7:0] out4704;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4704 = in0;
    end

    reg [7:0] out4705;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4705 = in0;
    end

    reg [7:0] out4706;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4706 = in0;
    end

    reg [7:0] out4707;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4707 = in0;
    end

    reg [7:0] out4708;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4708 = in0;
    end

    reg [7:0] out4709;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4709 = in0;
    end

    reg [7:0] out4710;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4710 = in0;
    end

    reg [7:0] out4711;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4711 = in0;
    end

    reg [7:0] out4712;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4712 = in0;
    end

    reg [7:0] out4713;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4713 = in0;
    end

    reg [7:0] out4714;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4714 = in0;
    end

    reg [7:0] out4715;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4715 = in0;
    end

    reg [7:0] out4716;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4716 = in0;
    end

    reg [7:0] out4717;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4717 = in0;
    end

    reg [7:0] out4718;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4718 = in0;
    end

    reg [7:0] out4719;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4719 = in0;
    end

    reg [7:0] out4720;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4720 = in0;
    end

    reg [7:0] out4721;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4721 = in0;
    end

    reg [7:0] out4722;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4722 = in0;
    end

    reg [7:0] out4723;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4723 = in0;
    end

    reg [7:0] out4724;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4724 = in0;
    end

    reg [7:0] out4725;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4725 = in0;
    end

    reg [7:0] out4726;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4726 = in0;
    end

    reg [7:0] out4727;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4727 = in0;
    end

    reg [7:0] out4728;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4728 = in0;
    end

    reg [7:0] out4729;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4729 = in0;
    end

    reg [7:0] out4730;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4730 = in0;
    end

    reg [7:0] out4731;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4731 = in0;
    end

    reg [7:0] out4732;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4732 = in0;
    end

    reg [7:0] out4733;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4733 = in0;
    end

    reg [7:0] out4734;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4734 = in0;
    end

    reg [7:0] out4735;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4735 = in0;
    end

    reg [7:0] out4736;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4736 = in0;
    end

    reg [7:0] out4737;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4737 = in0;
    end

    reg [7:0] out4738;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4738 = in0;
    end

    reg [7:0] out4739;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4739 = in0;
    end

    reg [7:0] out4740;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4740 = in0;
    end

    reg [7:0] out4741;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4741 = in0;
    end

    reg [7:0] out4742;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4742 = in0;
    end

    reg [7:0] out4743;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4743 = in0;
    end

    reg [7:0] out4744;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4744 = in0;
    end

    reg [7:0] out4745;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4745 = in0;
    end

    reg [7:0] out4746;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4746 = in0;
    end

    reg [7:0] out4747;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4747 = in0;
    end

    reg [7:0] out4748;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4748 = in0;
    end

    reg [7:0] out4749;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4749 = in0;
    end

    reg [7:0] out4750;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4750 = in0;
    end

    reg [7:0] out4751;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4751 = in0;
    end

    reg [7:0] out4752;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4752 = in0;
    end

    reg [7:0] out4753;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4753 = in0;
    end

    reg [7:0] out4754;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4754 = in0;
    end

    reg [7:0] out4755;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4755 = in0;
    end

    reg [7:0] out4756;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4756 = in0;
    end

    reg [7:0] out4757;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4757 = in0;
    end

    reg [7:0] out4758;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4758 = in0;
    end

    reg [7:0] out4759;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4759 = in0;
    end

    reg [7:0] out4760;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4760 = in0;
    end

    reg [7:0] out4761;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4761 = in0;
    end

    reg [7:0] out4762;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4762 = in0;
    end

    reg [7:0] out4763;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4763 = in0;
    end

    reg [7:0] out4764;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4764 = in0;
    end

    reg [7:0] out4765;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4765 = in0;
    end

    reg [7:0] out4766;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4766 = in0;
    end

    reg [7:0] out4767;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4767 = in0;
    end

    reg [7:0] out4768;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4768 = in0;
    end

    reg [7:0] out4769;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4769 = in0;
    end

    reg [7:0] out4770;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4770 = in0;
    end

    reg [7:0] out4771;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4771 = in0;
    end

    reg [7:0] out4772;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4772 = in0;
    end

    reg [7:0] out4773;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4773 = in0;
    end

    reg [7:0] out4774;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4774 = in0;
    end

    reg [7:0] out4775;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4775 = in0;
    end

    reg [7:0] out4776;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4776 = in0;
    end

    reg [7:0] out4777;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4777 = in0;
    end

    reg [7:0] out4778;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4778 = in0;
    end

    reg [7:0] out4779;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4779 = in0;
    end

    reg [7:0] out4780;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4780 = in0;
    end

    reg [7:0] out4781;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4781 = in0;
    end

    reg [7:0] out4782;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4782 = in0;
    end

    reg [7:0] out4783;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4783 = in0;
    end

    reg [7:0] out4784;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4784 = in0;
    end

    reg [7:0] out4785;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4785 = in0;
    end

    reg [7:0] out4786;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4786 = in0;
    end

    reg [7:0] out4787;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4787 = in0;
    end

    reg [7:0] out4788;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4788 = in0;
    end

    reg [7:0] out4789;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4789 = in0;
    end

    reg [7:0] out4790;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4790 = in0;
    end

    reg [7:0] out4791;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4791 = in0;
    end

    reg [7:0] out4792;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4792 = in0;
    end

    reg [7:0] out4793;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4793 = in0;
    end

    reg [7:0] out4794;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4794 = in0;
    end

    reg [7:0] out4795;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4795 = in0;
    end

    reg [7:0] out4796;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4796 = in0;
    end

    reg [7:0] out4797;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4797 = in0;
    end

    reg [7:0] out4798;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4798 = in0;
    end

    reg [7:0] out4799;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4799 = in0;
    end

    reg [7:0] out4800;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4800 = in0;
    end

    reg [7:0] out4801;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4801 = in0;
    end

    reg [7:0] out4802;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4802 = in0;
    end

    reg [7:0] out4803;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4803 = in0;
    end

    reg [7:0] out4804;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4804 = in0;
    end

    reg [7:0] out4805;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4805 = in0;
    end

    reg [7:0] out4806;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4806 = in0;
    end

    reg [7:0] out4807;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4807 = in0;
    end

    reg [7:0] out4808;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4808 = in0;
    end

    reg [7:0] out4809;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4809 = in0;
    end

    reg [7:0] out4810;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4810 = in0;
    end

    reg [7:0] out4811;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4811 = in0;
    end

    reg [7:0] out4812;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4812 = in0;
    end

    reg [7:0] out4813;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4813 = in0;
    end

    reg [7:0] out4814;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4814 = in0;
    end

    reg [7:0] out4815;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4815 = in0;
    end

    reg [7:0] out4816;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4816 = in0;
    end

    reg [7:0] out4817;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4817 = in0;
    end

    reg [7:0] out4818;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4818 = in0;
    end

    reg [7:0] out4819;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4819 = in0;
    end

    reg [7:0] out4820;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4820 = in0;
    end

    reg [7:0] out4821;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4821 = in0;
    end

    reg [7:0] out4822;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4822 = in0;
    end

    reg [7:0] out4823;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4823 = in0;
    end

    reg [7:0] out4824;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4824 = in0;
    end

    reg [7:0] out4825;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4825 = in0;
    end

    reg [7:0] out4826;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4826 = in0;
    end

    reg [7:0] out4827;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4827 = in0;
    end

    reg [7:0] out4828;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4828 = in0;
    end

    reg [7:0] out4829;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4829 = in0;
    end

    reg [7:0] out4830;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4830 = in0;
    end

    reg [7:0] out4831;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4831 = in0;
    end

    reg [7:0] out4832;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4832 = in0;
    end

    reg [7:0] out4833;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4833 = in0;
    end

    reg [7:0] out4834;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4834 = in0;
    end

    reg [7:0] out4835;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4835 = in0;
    end

    reg [7:0] out4836;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4836 = in0;
    end

    reg [7:0] out4837;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4837 = in0;
    end

    reg [7:0] out4838;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4838 = in0;
    end

    reg [7:0] out4839;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4839 = in0;
    end

    reg [7:0] out4840;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4840 = in0;
    end

    reg [7:0] out4841;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4841 = in0;
    end

    reg [7:0] out4842;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4842 = in0;
    end

    reg [7:0] out4843;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4843 = in0;
    end

    reg [7:0] out4844;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4844 = in0;
    end

    reg [7:0] out4845;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4845 = in0;
    end

    reg [7:0] out4846;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4846 = in0;
    end

    reg [7:0] out4847;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4847 = in0;
    end

    reg [7:0] out4848;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4848 = in0;
    end

    reg [7:0] out4849;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4849 = in0;
    end

    reg [7:0] out4850;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4850 = in0;
    end

    reg [7:0] out4851;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4851 = in0;
    end

    reg [7:0] out4852;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4852 = in0;
    end

    reg [7:0] out4853;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4853 = in0;
    end

    reg [7:0] out4854;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4854 = in0;
    end

    reg [7:0] out4855;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4855 = in0;
    end

    reg [7:0] out4856;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4856 = in0;
    end

    reg [7:0] out4857;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4857 = in0;
    end

    reg [7:0] out4858;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4858 = in0;
    end

    reg [7:0] out4859;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4859 = in0;
    end

    reg [7:0] out4860;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4860 = in0;
    end

    reg [7:0] out4861;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4861 = in0;
    end

    reg [7:0] out4862;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4862 = in0;
    end

    reg [7:0] out4863;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4863 = in0;
    end

    reg [7:0] out4864;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4864 = in0;
    end

    reg [7:0] out4865;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4865 = in0;
    end

    reg [7:0] out4866;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4866 = in0;
    end

    reg [7:0] out4867;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4867 = in0;
    end

    reg [7:0] out4868;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4868 = in0;
    end

    reg [7:0] out4869;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4869 = in0;
    end

    reg [7:0] out4870;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4870 = in0;
    end

    reg [7:0] out4871;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4871 = in0;
    end

    reg [7:0] out4872;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4872 = in0;
    end

    reg [7:0] out4873;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4873 = in0;
    end

    reg [7:0] out4874;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4874 = in0;
    end

    reg [7:0] out4875;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4875 = in0;
    end

    reg [7:0] out4876;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4876 = in0;
    end

    reg [7:0] out4877;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4877 = in0;
    end

    reg [7:0] out4878;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4878 = in0;
    end

    reg [7:0] out4879;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4879 = in0;
    end

    reg [7:0] out4880;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4880 = in0;
    end

    reg [7:0] out4881;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4881 = in0;
    end

    reg [7:0] out4882;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4882 = in0;
    end

    reg [7:0] out4883;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4883 = in0;
    end

    reg [7:0] out4884;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4884 = in0;
    end

    reg [7:0] out4885;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4885 = in0;
    end

    reg [7:0] out4886;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4886 = in0;
    end

    reg [7:0] out4887;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4887 = in0;
    end

    reg [7:0] out4888;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4888 = in0;
    end

    reg [7:0] out4889;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4889 = in0;
    end

    reg [7:0] out4890;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4890 = in0;
    end

    reg [7:0] out4891;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4891 = in0;
    end

    reg [7:0] out4892;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4892 = in0;
    end

    reg [7:0] out4893;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4893 = in0;
    end

    reg [7:0] out4894;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4894 = in0;
    end

    reg [7:0] out4895;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4895 = in0;
    end

    reg [7:0] out4896;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4896 = in0;
    end

    reg [7:0] out4897;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4897 = in0;
    end

    reg [7:0] out4898;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4898 = in0;
    end

    reg [7:0] out4899;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4899 = in0;
    end

    reg [7:0] out4900;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4900 = in0;
    end

    reg [7:0] out4901;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4901 = in0;
    end

    reg [7:0] out4902;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4902 = in0;
    end

    reg [7:0] out4903;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4903 = in0;
    end

    reg [7:0] out4904;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4904 = in0;
    end

    reg [7:0] out4905;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4905 = in0;
    end

    reg [7:0] out4906;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4906 = in0;
    end

    reg [7:0] out4907;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4907 = in0;
    end

    reg [7:0] out4908;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4908 = in0;
    end

    reg [7:0] out4909;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4909 = in0;
    end

    reg [7:0] out4910;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4910 = in0;
    end

    reg [7:0] out4911;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4911 = in0;
    end

    reg [7:0] out4912;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4912 = in0;
    end

    reg [7:0] out4913;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4913 = in0;
    end

    reg [7:0] out4914;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4914 = in0;
    end

    reg [7:0] out4915;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4915 = in0;
    end

    reg [7:0] out4916;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4916 = in0;
    end

    reg [7:0] out4917;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4917 = in0;
    end

    reg [7:0] out4918;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4918 = in0;
    end

    reg [7:0] out4919;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4919 = in0;
    end

    reg [7:0] out4920;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4920 = in0;
    end

    reg [7:0] out4921;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4921 = in0;
    end

    reg [7:0] out4922;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4922 = in0;
    end

    reg [7:0] out4923;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4923 = in0;
    end

    reg [7:0] out4924;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4924 = in0;
    end

    reg [7:0] out4925;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4925 = in0;
    end

    reg [7:0] out4926;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4926 = in0;
    end

    reg [7:0] out4927;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4927 = in0;
    end

    reg [7:0] out4928;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4928 = in0;
    end

    reg [7:0] out4929;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4929 = in0;
    end

    reg [7:0] out4930;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4930 = in0;
    end

    reg [7:0] out4931;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4931 = in0;
    end

    reg [7:0] out4932;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4932 = in0;
    end

    reg [7:0] out4933;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4933 = in0;
    end

    reg [7:0] out4934;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4934 = in0;
    end

    reg [7:0] out4935;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4935 = in0;
    end

    reg [7:0] out4936;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4936 = in0;
    end

    reg [7:0] out4937;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4937 = in0;
    end

    reg [7:0] out4938;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4938 = in0;
    end

    reg [7:0] out4939;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4939 = in0;
    end

    reg [7:0] out4940;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4940 = in0;
    end

    reg [7:0] out4941;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4941 = in0;
    end

    reg [7:0] out4942;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4942 = in0;
    end

    reg [7:0] out4943;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4943 = in0;
    end

    reg [7:0] out4944;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4944 = in0;
    end

    reg [7:0] out4945;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4945 = in0;
    end

    reg [7:0] out4946;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4946 = in0;
    end

    reg [7:0] out4947;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4947 = in0;
    end

    reg [7:0] out4948;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4948 = in0;
    end

    reg [7:0] out4949;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4949 = in0;
    end

    reg [7:0] out4950;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4950 = in0;
    end

    reg [7:0] out4951;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4951 = in0;
    end

    reg [7:0] out4952;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4952 = in0;
    end

    reg [7:0] out4953;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4953 = in0;
    end

    reg [7:0] out4954;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4954 = in0;
    end

    reg [7:0] out4955;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4955 = in0;
    end

    reg [7:0] out4956;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4956 = in0;
    end

    reg [7:0] out4957;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4957 = in0;
    end

    reg [7:0] out4958;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4958 = in0;
    end

    reg [7:0] out4959;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4959 = in0;
    end

    reg [7:0] out4960;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4960 = in0;
    end

    reg [7:0] out4961;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4961 = in0;
    end

    reg [7:0] out4962;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4962 = in0;
    end

    reg [7:0] out4963;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4963 = in0;
    end

    reg [7:0] out4964;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4964 = in0;
    end

    reg [7:0] out4965;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4965 = in0;
    end

    reg [7:0] out4966;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4966 = in0;
    end

    reg [7:0] out4967;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4967 = in0;
    end

    reg [7:0] out4968;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4968 = in0;
    end

    reg [7:0] out4969;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4969 = in0;
    end

    reg [7:0] out4970;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4970 = in0;
    end

    reg [7:0] out4971;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4971 = in0;
    end

    reg [7:0] out4972;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4972 = in0;
    end

    reg [7:0] out4973;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4973 = in0;
    end

    reg [7:0] out4974;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4974 = in0;
    end

    reg [7:0] out4975;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4975 = in0;
    end

    reg [7:0] out4976;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4976 = in0;
    end

    reg [7:0] out4977;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4977 = in0;
    end

    reg [7:0] out4978;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4978 = in0;
    end

    reg [7:0] out4979;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4979 = in0;
    end

    reg [7:0] out4980;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4980 = in0;
    end

    reg [7:0] out4981;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4981 = in0;
    end

    reg [7:0] out4982;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4982 = in0;
    end

    reg [7:0] out4983;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4983 = in0;
    end

    reg [7:0] out4984;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4984 = in0;
    end

    reg [7:0] out4985;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4985 = in0;
    end

    reg [7:0] out4986;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4986 = in0;
    end

    reg [7:0] out4987;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4987 = in0;
    end

    reg [7:0] out4988;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4988 = in0;
    end

    reg [7:0] out4989;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4989 = in0;
    end

    reg [7:0] out4990;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4990 = in0;
    end

    reg [7:0] out4991;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4991 = in0;
    end

    reg [7:0] out4992;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4992 = in0;
    end

    reg [7:0] out4993;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4993 = in0;
    end

    reg [7:0] out4994;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4994 = in0;
    end

    reg [7:0] out4995;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4995 = in0;
    end

    reg [7:0] out4996;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4996 = in0;
    end

    reg [7:0] out4997;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4997 = in0;
    end

    reg [7:0] out4998;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4998 = in0;
    end

    reg [7:0] out4999;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out4999 = in0;
    end

    reg [7:0] out5000;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5000 = in0;
    end

    reg [7:0] out5001;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5001 = in0;
    end

    reg [7:0] out5002;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5002 = in0;
    end

    reg [7:0] out5003;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5003 = in0;
    end

    reg [7:0] out5004;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5004 = in0;
    end

    reg [7:0] out5005;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5005 = in0;
    end

    reg [7:0] out5006;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5006 = in0;
    end

    reg [7:0] out5007;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5007 = in0;
    end

    reg [7:0] out5008;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5008 = in0;
    end

    reg [7:0] out5009;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5009 = in0;
    end

    reg [7:0] out5010;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5010 = in0;
    end

    reg [7:0] out5011;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5011 = in0;
    end

    reg [7:0] out5012;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5012 = in0;
    end

    reg [7:0] out5013;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5013 = in0;
    end

    reg [7:0] out5014;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5014 = in0;
    end

    reg [7:0] out5015;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5015 = in0;
    end

    reg [7:0] out5016;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5016 = in0;
    end

    reg [7:0] out5017;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5017 = in0;
    end

    reg [7:0] out5018;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5018 = in0;
    end

    reg [7:0] out5019;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5019 = in0;
    end

    reg [7:0] out5020;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5020 = in0;
    end

    reg [7:0] out5021;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5021 = in0;
    end

    reg [7:0] out5022;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5022 = in0;
    end

    reg [7:0] out5023;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5023 = in0;
    end

    reg [7:0] out5024;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5024 = in0;
    end

    reg [7:0] out5025;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5025 = in0;
    end

    reg [7:0] out5026;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5026 = in0;
    end

    reg [7:0] out5027;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5027 = in0;
    end

    reg [7:0] out5028;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5028 = in0;
    end

    reg [7:0] out5029;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5029 = in0;
    end

    reg [7:0] out5030;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5030 = in0;
    end

    reg [7:0] out5031;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5031 = in0;
    end

    reg [7:0] out5032;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5032 = in0;
    end

    reg [7:0] out5033;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5033 = in0;
    end

    reg [7:0] out5034;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5034 = in0;
    end

    reg [7:0] out5035;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5035 = in0;
    end

    reg [7:0] out5036;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5036 = in0;
    end

    reg [7:0] out5037;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5037 = in0;
    end

    reg [7:0] out5038;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5038 = in0;
    end

    reg [7:0] out5039;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5039 = in0;
    end

    reg [7:0] out5040;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5040 = in0;
    end

    reg [7:0] out5041;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5041 = in0;
    end

    reg [7:0] out5042;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5042 = in0;
    end

    reg [7:0] out5043;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5043 = in0;
    end

    reg [7:0] out5044;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5044 = in0;
    end

    reg [7:0] out5045;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5045 = in0;
    end

    reg [7:0] out5046;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5046 = in0;
    end

    reg [7:0] out5047;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5047 = in0;
    end

    reg [7:0] out5048;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5048 = in0;
    end

    reg [7:0] out5049;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5049 = in0;
    end

    reg [7:0] out5050;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5050 = in0;
    end

    reg [7:0] out5051;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5051 = in0;
    end

    reg [7:0] out5052;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5052 = in0;
    end

    reg [7:0] out5053;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5053 = in0;
    end

    reg [7:0] out5054;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5054 = in0;
    end

    reg [7:0] out5055;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5055 = in0;
    end

    reg [7:0] out5056;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5056 = in0;
    end

    reg [7:0] out5057;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5057 = in0;
    end

    reg [7:0] out5058;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5058 = in0;
    end

    reg [7:0] out5059;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5059 = in0;
    end

    reg [7:0] out5060;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5060 = in0;
    end

    reg [7:0] out5061;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5061 = in0;
    end

    reg [7:0] out5062;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5062 = in0;
    end

    reg [7:0] out5063;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5063 = in0;
    end

    reg [7:0] out5064;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5064 = in0;
    end

    reg [7:0] out5065;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5065 = in0;
    end

    reg [7:0] out5066;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5066 = in0;
    end

    reg [7:0] out5067;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5067 = in0;
    end

    reg [7:0] out5068;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5068 = in0;
    end

    reg [7:0] out5069;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5069 = in0;
    end

    reg [7:0] out5070;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5070 = in0;
    end

    reg [7:0] out5071;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5071 = in0;
    end

    reg [7:0] out5072;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5072 = in0;
    end

    reg [7:0] out5073;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5073 = in0;
    end

    reg [7:0] out5074;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5074 = in0;
    end

    reg [7:0] out5075;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5075 = in0;
    end

    reg [7:0] out5076;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5076 = in0;
    end

    reg [7:0] out5077;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5077 = in0;
    end

    reg [7:0] out5078;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5078 = in0;
    end

    reg [7:0] out5079;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5079 = in0;
    end

    reg [7:0] out5080;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5080 = in0;
    end

    reg [7:0] out5081;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5081 = in0;
    end

    reg [7:0] out5082;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5082 = in0;
    end

    reg [7:0] out5083;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5083 = in0;
    end

    reg [7:0] out5084;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5084 = in0;
    end

    reg [7:0] out5085;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5085 = in0;
    end

    reg [7:0] out5086;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5086 = in0;
    end

    reg [7:0] out5087;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5087 = in0;
    end

    reg [7:0] out5088;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5088 = in0;
    end

    reg [7:0] out5089;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5089 = in0;
    end

    reg [7:0] out5090;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5090 = in0;
    end

    reg [7:0] out5091;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5091 = in0;
    end

    reg [7:0] out5092;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5092 = in0;
    end

    reg [7:0] out5093;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5093 = in0;
    end

    reg [7:0] out5094;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5094 = in0;
    end

    reg [7:0] out5095;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5095 = in0;
    end

    reg [7:0] out5096;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5096 = in0;
    end

    reg [7:0] out5097;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5097 = in0;
    end

    reg [7:0] out5098;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5098 = in0;
    end

    reg [7:0] out5099;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5099 = in0;
    end

    reg [7:0] out5100;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5100 = in0;
    end

    reg [7:0] out5101;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5101 = in0;
    end

    reg [7:0] out5102;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5102 = in0;
    end

    reg [7:0] out5103;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5103 = in0;
    end

    reg [7:0] out5104;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5104 = in0;
    end

    reg [7:0] out5105;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5105 = in0;
    end

    reg [7:0] out5106;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5106 = in0;
    end

    reg [7:0] out5107;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5107 = in0;
    end

    reg [7:0] out5108;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5108 = in0;
    end

    reg [7:0] out5109;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5109 = in0;
    end

    reg [7:0] out5110;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5110 = in0;
    end

    reg [7:0] out5111;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5111 = in0;
    end

    reg [7:0] out5112;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5112 = in0;
    end

    reg [7:0] out5113;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5113 = in0;
    end

    reg [7:0] out5114;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5114 = in0;
    end

    reg [7:0] out5115;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5115 = in0;
    end

    reg [7:0] out5116;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5116 = in0;
    end

    reg [7:0] out5117;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5117 = in0;
    end

    reg [7:0] out5118;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5118 = in0;
    end

    reg [7:0] out5119;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5119 = in0;
    end

    reg [7:0] out5120;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5120 = in0;
    end

    reg [7:0] out5121;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5121 = in0;
    end

    reg [7:0] out5122;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5122 = in0;
    end

    reg [7:0] out5123;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5123 = in0;
    end

    reg [7:0] out5124;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5124 = in0;
    end

    reg [7:0] out5125;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5125 = in0;
    end

    reg [7:0] out5126;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5126 = in0;
    end

    reg [7:0] out5127;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5127 = in0;
    end

    reg [7:0] out5128;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5128 = in0;
    end

    reg [7:0] out5129;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5129 = in0;
    end

    reg [7:0] out5130;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5130 = in0;
    end

    reg [7:0] out5131;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5131 = in0;
    end

    reg [7:0] out5132;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5132 = in0;
    end

    reg [7:0] out5133;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5133 = in0;
    end

    reg [7:0] out5134;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5134 = in0;
    end

    reg [7:0] out5135;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5135 = in0;
    end

    reg [7:0] out5136;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5136 = in0;
    end

    reg [7:0] out5137;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5137 = in0;
    end

    reg [7:0] out5138;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5138 = in0;
    end

    reg [7:0] out5139;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5139 = in0;
    end

    reg [7:0] out5140;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5140 = in0;
    end

    reg [7:0] out5141;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5141 = in0;
    end

    reg [7:0] out5142;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5142 = in0;
    end

    reg [7:0] out5143;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5143 = in0;
    end

    reg [7:0] out5144;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5144 = in0;
    end

    reg [7:0] out5145;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5145 = in0;
    end

    reg [7:0] out5146;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5146 = in0;
    end

    reg [7:0] out5147;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5147 = in0;
    end

    reg [7:0] out5148;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5148 = in0;
    end

    reg [7:0] out5149;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5149 = in0;
    end

    reg [7:0] out5150;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5150 = in0;
    end

    reg [7:0] out5151;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5151 = in0;
    end

    reg [7:0] out5152;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5152 = in0;
    end

    reg [7:0] out5153;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5153 = in0;
    end

    reg [7:0] out5154;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5154 = in0;
    end

    reg [7:0] out5155;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5155 = in0;
    end

    reg [7:0] out5156;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5156 = in0;
    end

    reg [7:0] out5157;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5157 = in0;
    end

    reg [7:0] out5158;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5158 = in0;
    end

    reg [7:0] out5159;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5159 = in0;
    end

    reg [7:0] out5160;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5160 = in0;
    end

    reg [7:0] out5161;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5161 = in0;
    end

    reg [7:0] out5162;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5162 = in0;
    end

    reg [7:0] out5163;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5163 = in0;
    end

    reg [7:0] out5164;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5164 = in0;
    end

    reg [7:0] out5165;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5165 = in0;
    end

    reg [7:0] out5166;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5166 = in0;
    end

    reg [7:0] out5167;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5167 = in0;
    end

    reg [7:0] out5168;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5168 = in0;
    end

    reg [7:0] out5169;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5169 = in0;
    end

    reg [7:0] out5170;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5170 = in0;
    end

    reg [7:0] out5171;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5171 = in0;
    end

    reg [7:0] out5172;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5172 = in0;
    end

    reg [7:0] out5173;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5173 = in0;
    end

    reg [7:0] out5174;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5174 = in0;
    end

    reg [7:0] out5175;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5175 = in0;
    end

    reg [7:0] out5176;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5176 = in0;
    end

    reg [7:0] out5177;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5177 = in0;
    end

    reg [7:0] out5178;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5178 = in0;
    end

    reg [7:0] out5179;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5179 = in0;
    end

    reg [7:0] out5180;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5180 = in0;
    end

    reg [7:0] out5181;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5181 = in0;
    end

    reg [7:0] out5182;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5182 = in0;
    end

    reg [7:0] out5183;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5183 = in0;
    end

    reg [7:0] out5184;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5184 = in0;
    end

    reg [7:0] out5185;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5185 = in0;
    end

    reg [7:0] out5186;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5186 = in0;
    end

    reg [7:0] out5187;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5187 = in0;
    end

    reg [7:0] out5188;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5188 = in0;
    end

    reg [7:0] out5189;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5189 = in0;
    end

    reg [7:0] out5190;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5190 = in0;
    end

    reg [7:0] out5191;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5191 = in0;
    end

    reg [7:0] out5192;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5192 = in0;
    end

    reg [7:0] out5193;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5193 = in0;
    end

    reg [7:0] out5194;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5194 = in0;
    end

    reg [7:0] out5195;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5195 = in0;
    end

    reg [7:0] out5196;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5196 = in0;
    end

    reg [7:0] out5197;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5197 = in0;
    end

    reg [7:0] out5198;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5198 = in0;
    end

    reg [7:0] out5199;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5199 = in0;
    end

    reg [7:0] out5200;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5200 = in0;
    end

    reg [7:0] out5201;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5201 = in0;
    end

    reg [7:0] out5202;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5202 = in0;
    end

    reg [7:0] out5203;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5203 = in0;
    end

    reg [7:0] out5204;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5204 = in0;
    end

    reg [7:0] out5205;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5205 = in0;
    end

    reg [7:0] out5206;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5206 = in0;
    end

    reg [7:0] out5207;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5207 = in0;
    end

    reg [7:0] out5208;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5208 = in0;
    end

    reg [7:0] out5209;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5209 = in0;
    end

    reg [7:0] out5210;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5210 = in0;
    end

    reg [7:0] out5211;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5211 = in0;
    end

    reg [7:0] out5212;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5212 = in0;
    end

    reg [7:0] out5213;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5213 = in0;
    end

    reg [7:0] out5214;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5214 = in0;
    end

    reg [7:0] out5215;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5215 = in0;
    end

    reg [7:0] out5216;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5216 = in0;
    end

    reg [7:0] out5217;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5217 = in0;
    end

    reg [7:0] out5218;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5218 = in0;
    end

    reg [7:0] out5219;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5219 = in0;
    end

    reg [7:0] out5220;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5220 = in0;
    end

    reg [7:0] out5221;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5221 = in0;
    end

    reg [7:0] out5222;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5222 = in0;
    end

    reg [7:0] out5223;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5223 = in0;
    end

    reg [7:0] out5224;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5224 = in0;
    end

    reg [7:0] out5225;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5225 = in0;
    end

    reg [7:0] out5226;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5226 = in0;
    end

    reg [7:0] out5227;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5227 = in0;
    end

    reg [7:0] out5228;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5228 = in0;
    end

    reg [7:0] out5229;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5229 = in0;
    end

    reg [7:0] out5230;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5230 = in0;
    end

    reg [7:0] out5231;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5231 = in0;
    end

    reg [7:0] out5232;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5232 = in0;
    end

    reg [7:0] out5233;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5233 = in0;
    end

    reg [7:0] out5234;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5234 = in0;
    end

    reg [7:0] out5235;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5235 = in0;
    end

    reg [7:0] out5236;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5236 = in0;
    end

    reg [7:0] out5237;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5237 = in0;
    end

    reg [7:0] out5238;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5238 = in0;
    end

    reg [7:0] out5239;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5239 = in0;
    end

    reg [7:0] out5240;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5240 = in0;
    end

    reg [7:0] out5241;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5241 = in0;
    end

    reg [7:0] out5242;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5242 = in0;
    end

    reg [7:0] out5243;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5243 = in0;
    end

    reg [7:0] out5244;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5244 = in0;
    end

    reg [7:0] out5245;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5245 = in0;
    end

    reg [7:0] out5246;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5246 = in0;
    end

    reg [7:0] out5247;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5247 = in0;
    end

    reg [7:0] out5248;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5248 = in0;
    end

    reg [7:0] out5249;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5249 = in0;
    end

    reg [7:0] out5250;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5250 = in0;
    end

    reg [7:0] out5251;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5251 = in0;
    end

    reg [7:0] out5252;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5252 = in0;
    end

    reg [7:0] out5253;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5253 = in0;
    end

    reg [7:0] out5254;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5254 = in0;
    end

    reg [7:0] out5255;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5255 = in0;
    end

    reg [7:0] out5256;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5256 = in0;
    end

    reg [7:0] out5257;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5257 = in0;
    end

    reg [7:0] out5258;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5258 = in0;
    end

    reg [7:0] out5259;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5259 = in0;
    end

    reg [7:0] out5260;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5260 = in0;
    end

    reg [7:0] out5261;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5261 = in0;
    end

    reg [7:0] out5262;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5262 = in0;
    end

    reg [7:0] out5263;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5263 = in0;
    end

    reg [7:0] out5264;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5264 = in0;
    end

    reg [7:0] out5265;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5265 = in0;
    end

    reg [7:0] out5266;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5266 = in0;
    end

    reg [7:0] out5267;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5267 = in0;
    end

    reg [7:0] out5268;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5268 = in0;
    end

    reg [7:0] out5269;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5269 = in0;
    end

    reg [7:0] out5270;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5270 = in0;
    end

    reg [7:0] out5271;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5271 = in0;
    end

    reg [7:0] out5272;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5272 = in0;
    end

    reg [7:0] out5273;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5273 = in0;
    end

    reg [7:0] out5274;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5274 = in0;
    end

    reg [7:0] out5275;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5275 = in0;
    end

    reg [7:0] out5276;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5276 = in0;
    end

    reg [7:0] out5277;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5277 = in0;
    end

    reg [7:0] out5278;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5278 = in0;
    end

    reg [7:0] out5279;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5279 = in0;
    end

    reg [7:0] out5280;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5280 = in0;
    end

    reg [7:0] out5281;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5281 = in0;
    end

    reg [7:0] out5282;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5282 = in0;
    end

    reg [7:0] out5283;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5283 = in0;
    end

    reg [7:0] out5284;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5284 = in0;
    end

    reg [7:0] out5285;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5285 = in0;
    end

    reg [7:0] out5286;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5286 = in0;
    end

    reg [7:0] out5287;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5287 = in0;
    end

    reg [7:0] out5288;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5288 = in0;
    end

    reg [7:0] out5289;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5289 = in0;
    end

    reg [7:0] out5290;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5290 = in0;
    end

    reg [7:0] out5291;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5291 = in0;
    end

    reg [7:0] out5292;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5292 = in0;
    end

    reg [7:0] out5293;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5293 = in0;
    end

    reg [7:0] out5294;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5294 = in0;
    end

    reg [7:0] out5295;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5295 = in0;
    end

    reg [7:0] out5296;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5296 = in0;
    end

    reg [7:0] out5297;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5297 = in0;
    end

    reg [7:0] out5298;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5298 = in0;
    end

    reg [7:0] out5299;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5299 = in0;
    end

    reg [7:0] out5300;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5300 = in0;
    end

    reg [7:0] out5301;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5301 = in0;
    end

    reg [7:0] out5302;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5302 = in0;
    end

    reg [7:0] out5303;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5303 = in0;
    end

    reg [7:0] out5304;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5304 = in0;
    end

    reg [7:0] out5305;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5305 = in0;
    end

    reg [7:0] out5306;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5306 = in0;
    end

    reg [7:0] out5307;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5307 = in0;
    end

    reg [7:0] out5308;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5308 = in0;
    end

    reg [7:0] out5309;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5309 = in0;
    end

    reg [7:0] out5310;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5310 = in0;
    end

    reg [7:0] out5311;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5311 = in0;
    end

    reg [7:0] out5312;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5312 = in0;
    end

    reg [7:0] out5313;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5313 = in0;
    end

    reg [7:0] out5314;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5314 = in0;
    end

    reg [7:0] out5315;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5315 = in0;
    end

    reg [7:0] out5316;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5316 = in0;
    end

    reg [7:0] out5317;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5317 = in0;
    end

    reg [7:0] out5318;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5318 = in0;
    end

    reg [7:0] out5319;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5319 = in0;
    end

    reg [7:0] out5320;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5320 = in0;
    end

    reg [7:0] out5321;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5321 = in0;
    end

    reg [7:0] out5322;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5322 = in0;
    end

    reg [7:0] out5323;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5323 = in0;
    end

    reg [7:0] out5324;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5324 = in0;
    end

    reg [7:0] out5325;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5325 = in0;
    end

    reg [7:0] out5326;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5326 = in0;
    end

    reg [7:0] out5327;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5327 = in0;
    end

    reg [7:0] out5328;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5328 = in0;
    end

    reg [7:0] out5329;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5329 = in0;
    end

    reg [7:0] out5330;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5330 = in0;
    end

    reg [7:0] out5331;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5331 = in0;
    end

    reg [7:0] out5332;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5332 = in0;
    end

    reg [7:0] out5333;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5333 = in0;
    end

    reg [7:0] out5334;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5334 = in0;
    end

    reg [7:0] out5335;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5335 = in0;
    end

    reg [7:0] out5336;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5336 = in0;
    end

    reg [7:0] out5337;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5337 = in0;
    end

    reg [7:0] out5338;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5338 = in0;
    end

    reg [7:0] out5339;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5339 = in0;
    end

    reg [7:0] out5340;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5340 = in0;
    end

    reg [7:0] out5341;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5341 = in0;
    end

    reg [7:0] out5342;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5342 = in0;
    end

    reg [7:0] out5343;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5343 = in0;
    end

    reg [7:0] out5344;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5344 = in0;
    end

    reg [7:0] out5345;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5345 = in0;
    end

    reg [7:0] out5346;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5346 = in0;
    end

    reg [7:0] out5347;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5347 = in0;
    end

    reg [7:0] out5348;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5348 = in0;
    end

    reg [7:0] out5349;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5349 = in0;
    end

    reg [7:0] out5350;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5350 = in0;
    end

    reg [7:0] out5351;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5351 = in0;
    end

    reg [7:0] out5352;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5352 = in0;
    end

    reg [7:0] out5353;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5353 = in0;
    end

    reg [7:0] out5354;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5354 = in0;
    end

    reg [7:0] out5355;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5355 = in0;
    end

    reg [7:0] out5356;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5356 = in0;
    end

    reg [7:0] out5357;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5357 = in0;
    end

    reg [7:0] out5358;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5358 = in0;
    end

    reg [7:0] out5359;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5359 = in0;
    end

    reg [7:0] out5360;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5360 = in0;
    end

    reg [7:0] out5361;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5361 = in0;
    end

    reg [7:0] out5362;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5362 = in0;
    end

    reg [7:0] out5363;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5363 = in0;
    end

    reg [7:0] out5364;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5364 = in0;
    end

    reg [7:0] out5365;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5365 = in0;
    end

    reg [7:0] out5366;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5366 = in0;
    end

    reg [7:0] out5367;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5367 = in0;
    end

    reg [7:0] out5368;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5368 = in0;
    end

    reg [7:0] out5369;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5369 = in0;
    end

    reg [7:0] out5370;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5370 = in0;
    end

    reg [7:0] out5371;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5371 = in0;
    end

    reg [7:0] out5372;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5372 = in0;
    end

    reg [7:0] out5373;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5373 = in0;
    end

    reg [7:0] out5374;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5374 = in0;
    end

    reg [7:0] out5375;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5375 = in0;
    end

    reg [7:0] out5376;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5376 = in0;
    end

    reg [7:0] out5377;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5377 = in0;
    end

    reg [7:0] out5378;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5378 = in0;
    end

    reg [7:0] out5379;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5379 = in0;
    end

    reg [7:0] out5380;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5380 = in0;
    end

    reg [7:0] out5381;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5381 = in0;
    end

    reg [7:0] out5382;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5382 = in0;
    end

    reg [7:0] out5383;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5383 = in0;
    end

    reg [7:0] out5384;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5384 = in0;
    end

    reg [7:0] out5385;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5385 = in0;
    end

    reg [7:0] out5386;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5386 = in0;
    end

    reg [7:0] out5387;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5387 = in0;
    end

    reg [7:0] out5388;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5388 = in0;
    end

    reg [7:0] out5389;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5389 = in0;
    end

    reg [7:0] out5390;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5390 = in0;
    end

    reg [7:0] out5391;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5391 = in0;
    end

    reg [7:0] out5392;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5392 = in0;
    end

    reg [7:0] out5393;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5393 = in0;
    end

    reg [7:0] out5394;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5394 = in0;
    end

    reg [7:0] out5395;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5395 = in0;
    end

    reg [7:0] out5396;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5396 = in0;
    end

    reg [7:0] out5397;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5397 = in0;
    end

    reg [7:0] out5398;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5398 = in0;
    end

    reg [7:0] out5399;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5399 = in0;
    end

    reg [7:0] out5400;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5400 = in0;
    end

    reg [7:0] out5401;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5401 = in0;
    end

    reg [7:0] out5402;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5402 = in0;
    end

    reg [7:0] out5403;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5403 = in0;
    end

    reg [7:0] out5404;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5404 = in0;
    end

    reg [7:0] out5405;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5405 = in0;
    end

    reg [7:0] out5406;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5406 = in0;
    end

    reg [7:0] out5407;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5407 = in0;
    end

    reg [7:0] out5408;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5408 = in0;
    end

    reg [7:0] out5409;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5409 = in0;
    end

    reg [7:0] out5410;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5410 = in0;
    end

    reg [7:0] out5411;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5411 = in0;
    end

    reg [7:0] out5412;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5412 = in0;
    end

    reg [7:0] out5413;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5413 = in0;
    end

    reg [7:0] out5414;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5414 = in0;
    end

    reg [7:0] out5415;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5415 = in0;
    end

    reg [7:0] out5416;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5416 = in0;
    end

    reg [7:0] out5417;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5417 = in0;
    end

    reg [7:0] out5418;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5418 = in0;
    end

    reg [7:0] out5419;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5419 = in0;
    end

    reg [7:0] out5420;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5420 = in0;
    end

    reg [7:0] out5421;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5421 = in0;
    end

    reg [7:0] out5422;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5422 = in0;
    end

    reg [7:0] out5423;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5423 = in0;
    end

    reg [7:0] out5424;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5424 = in0;
    end

    reg [7:0] out5425;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5425 = in0;
    end

    reg [7:0] out5426;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5426 = in0;
    end

    reg [7:0] out5427;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5427 = in0;
    end

    reg [7:0] out5428;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5428 = in0;
    end

    reg [7:0] out5429;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5429 = in0;
    end

    reg [7:0] out5430;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5430 = in0;
    end

    reg [7:0] out5431;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5431 = in0;
    end

    reg [7:0] out5432;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5432 = in0;
    end

    reg [7:0] out5433;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5433 = in0;
    end

    reg [7:0] out5434;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5434 = in0;
    end

    reg [7:0] out5435;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5435 = in0;
    end

    reg [7:0] out5436;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5436 = in0;
    end

    reg [7:0] out5437;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5437 = in0;
    end

    reg [7:0] out5438;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5438 = in0;
    end

    reg [7:0] out5439;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5439 = in0;
    end

    reg [7:0] out5440;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5440 = in0;
    end

    reg [7:0] out5441;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5441 = in0;
    end

    reg [7:0] out5442;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5442 = in0;
    end

    reg [7:0] out5443;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5443 = in0;
    end

    reg [7:0] out5444;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5444 = in0;
    end

    reg [7:0] out5445;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5445 = in0;
    end

    reg [7:0] out5446;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5446 = in0;
    end

    reg [7:0] out5447;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5447 = in0;
    end

    reg [7:0] out5448;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5448 = in0;
    end

    reg [7:0] out5449;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5449 = in0;
    end

    reg [7:0] out5450;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5450 = in0;
    end

    reg [7:0] out5451;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5451 = in0;
    end

    reg [7:0] out5452;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5452 = in0;
    end

    reg [7:0] out5453;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5453 = in0;
    end

    reg [7:0] out5454;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5454 = in0;
    end

    reg [7:0] out5455;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5455 = in0;
    end

    reg [7:0] out5456;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5456 = in0;
    end

    reg [7:0] out5457;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5457 = in0;
    end

    reg [7:0] out5458;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5458 = in0;
    end

    reg [7:0] out5459;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5459 = in0;
    end

    reg [7:0] out5460;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5460 = in0;
    end

    reg [7:0] out5461;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5461 = in0;
    end

    reg [7:0] out5462;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5462 = in0;
    end

    reg [7:0] out5463;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5463 = in0;
    end

    reg [7:0] out5464;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5464 = in0;
    end

    reg [7:0] out5465;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5465 = in0;
    end

    reg [7:0] out5466;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5466 = in0;
    end

    reg [7:0] out5467;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5467 = in0;
    end

    reg [7:0] out5468;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5468 = in0;
    end

    reg [7:0] out5469;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5469 = in0;
    end

    reg [7:0] out5470;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5470 = in0;
    end

    reg [7:0] out5471;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5471 = in0;
    end

    reg [7:0] out5472;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5472 = in0;
    end

    reg [7:0] out5473;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5473 = in0;
    end

    reg [7:0] out5474;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5474 = in0;
    end

    reg [7:0] out5475;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5475 = in0;
    end

    reg [7:0] out5476;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5476 = in0;
    end

    reg [7:0] out5477;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5477 = in0;
    end

    reg [7:0] out5478;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5478 = in0;
    end

    reg [7:0] out5479;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5479 = in0;
    end

    reg [7:0] out5480;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5480 = in0;
    end

    reg [7:0] out5481;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5481 = in0;
    end

    reg [7:0] out5482;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5482 = in0;
    end

    reg [7:0] out5483;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5483 = in0;
    end

    reg [7:0] out5484;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5484 = in0;
    end

    reg [7:0] out5485;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5485 = in0;
    end

    reg [7:0] out5486;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5486 = in0;
    end

    reg [7:0] out5487;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5487 = in0;
    end

    reg [7:0] out5488;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5488 = in0;
    end

    reg [7:0] out5489;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5489 = in0;
    end

    reg [7:0] out5490;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5490 = in0;
    end

    reg [7:0] out5491;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5491 = in0;
    end

    reg [7:0] out5492;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5492 = in0;
    end

    reg [7:0] out5493;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5493 = in0;
    end

    reg [7:0] out5494;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5494 = in0;
    end

    reg [7:0] out5495;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5495 = in0;
    end

    reg [7:0] out5496;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5496 = in0;
    end

    reg [7:0] out5497;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5497 = in0;
    end

    reg [7:0] out5498;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5498 = in0;
    end

    reg [7:0] out5499;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5499 = in0;
    end

    reg [7:0] out5500;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5500 = in0;
    end

    reg [7:0] out5501;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5501 = in0;
    end

    reg [7:0] out5502;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5502 = in0;
    end

    reg [7:0] out5503;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5503 = in0;
    end

    reg [7:0] out5504;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5504 = in0;
    end

    reg [7:0] out5505;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5505 = in0;
    end

    reg [7:0] out5506;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5506 = in0;
    end

    reg [7:0] out5507;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5507 = in0;
    end

    reg [7:0] out5508;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5508 = in0;
    end

    reg [7:0] out5509;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5509 = in0;
    end

    reg [7:0] out5510;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5510 = in0;
    end

    reg [7:0] out5511;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5511 = in0;
    end

    reg [7:0] out5512;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5512 = in0;
    end

    reg [7:0] out5513;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5513 = in0;
    end

    reg [7:0] out5514;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5514 = in0;
    end

    reg [7:0] out5515;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5515 = in0;
    end

    reg [7:0] out5516;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5516 = in0;
    end

    reg [7:0] out5517;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5517 = in0;
    end

    reg [7:0] out5518;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5518 = in0;
    end

    reg [7:0] out5519;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5519 = in0;
    end

    reg [7:0] out5520;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5520 = in0;
    end

    reg [7:0] out5521;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5521 = in0;
    end

    reg [7:0] out5522;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5522 = in0;
    end

    reg [7:0] out5523;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5523 = in0;
    end

    reg [7:0] out5524;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5524 = in0;
    end

    reg [7:0] out5525;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5525 = in0;
    end

    reg [7:0] out5526;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5526 = in0;
    end

    reg [7:0] out5527;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5527 = in0;
    end

    reg [7:0] out5528;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5528 = in0;
    end

    reg [7:0] out5529;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5529 = in0;
    end

    reg [7:0] out5530;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5530 = in0;
    end

    reg [7:0] out5531;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5531 = in0;
    end

    reg [7:0] out5532;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5532 = in0;
    end

    reg [7:0] out5533;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5533 = in0;
    end

    reg [7:0] out5534;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5534 = in0;
    end

    reg [7:0] out5535;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5535 = in0;
    end

    reg [7:0] out5536;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5536 = in0;
    end

    reg [7:0] out5537;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5537 = in0;
    end

    reg [7:0] out5538;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5538 = in0;
    end

    reg [7:0] out5539;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5539 = in0;
    end

    reg [7:0] out5540;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5540 = in0;
    end

    reg [7:0] out5541;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5541 = in0;
    end

    reg [7:0] out5542;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5542 = in0;
    end

    reg [7:0] out5543;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5543 = in0;
    end

    reg [7:0] out5544;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5544 = in0;
    end

    reg [7:0] out5545;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5545 = in0;
    end

    reg [7:0] out5546;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5546 = in0;
    end

    reg [7:0] out5547;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5547 = in0;
    end

    reg [7:0] out5548;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5548 = in0;
    end

    reg [7:0] out5549;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5549 = in0;
    end

    reg [7:0] out5550;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5550 = in0;
    end

    reg [7:0] out5551;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5551 = in0;
    end

    reg [7:0] out5552;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5552 = in0;
    end

    reg [7:0] out5553;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5553 = in0;
    end

    reg [7:0] out5554;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5554 = in0;
    end

    reg [7:0] out5555;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5555 = in0;
    end

    reg [7:0] out5556;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5556 = in0;
    end

    reg [7:0] out5557;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5557 = in0;
    end

    reg [7:0] out5558;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5558 = in0;
    end

    reg [7:0] out5559;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5559 = in0;
    end

    reg [7:0] out5560;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5560 = in0;
    end

    reg [7:0] out5561;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5561 = in0;
    end

    reg [7:0] out5562;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5562 = in0;
    end

    reg [7:0] out5563;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5563 = in0;
    end

    reg [7:0] out5564;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5564 = in0;
    end

    reg [7:0] out5565;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5565 = in0;
    end

    reg [7:0] out5566;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5566 = in0;
    end

    reg [7:0] out5567;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5567 = in0;
    end

    reg [7:0] out5568;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5568 = in0;
    end

    reg [7:0] out5569;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5569 = in0;
    end

    reg [7:0] out5570;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5570 = in0;
    end

    reg [7:0] out5571;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5571 = in0;
    end

    reg [7:0] out5572;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5572 = in0;
    end

    reg [7:0] out5573;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5573 = in0;
    end

    reg [7:0] out5574;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5574 = in0;
    end

    reg [7:0] out5575;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5575 = in0;
    end

    reg [7:0] out5576;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5576 = in0;
    end

    reg [7:0] out5577;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5577 = in0;
    end

    reg [7:0] out5578;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5578 = in0;
    end

    reg [7:0] out5579;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5579 = in0;
    end

    reg [7:0] out5580;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5580 = in0;
    end

    reg [7:0] out5581;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5581 = in0;
    end

    reg [7:0] out5582;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5582 = in0;
    end

    reg [7:0] out5583;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5583 = in0;
    end

    reg [7:0] out5584;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5584 = in0;
    end

    reg [7:0] out5585;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5585 = in0;
    end

    reg [7:0] out5586;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5586 = in0;
    end

    reg [7:0] out5587;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5587 = in0;
    end

    reg [7:0] out5588;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5588 = in0;
    end

    reg [7:0] out5589;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5589 = in0;
    end

    reg [7:0] out5590;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5590 = in0;
    end

    reg [7:0] out5591;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5591 = in0;
    end

    reg [7:0] out5592;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5592 = in0;
    end

    reg [7:0] out5593;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5593 = in0;
    end

    reg [7:0] out5594;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5594 = in0;
    end

    reg [7:0] out5595;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5595 = in0;
    end

    reg [7:0] out5596;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5596 = in0;
    end

    reg [7:0] out5597;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5597 = in0;
    end

    reg [7:0] out5598;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5598 = in0;
    end

    reg [7:0] out5599;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5599 = in0;
    end

    reg [7:0] out5600;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5600 = in0;
    end

    reg [7:0] out5601;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5601 = in0;
    end

    reg [7:0] out5602;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5602 = in0;
    end

    reg [7:0] out5603;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5603 = in0;
    end

    reg [7:0] out5604;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5604 = in0;
    end

    reg [7:0] out5605;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5605 = in0;
    end

    reg [7:0] out5606;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5606 = in0;
    end

    reg [7:0] out5607;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5607 = in0;
    end

    reg [7:0] out5608;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5608 = in0;
    end

    reg [7:0] out5609;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5609 = in0;
    end

    reg [7:0] out5610;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5610 = in0;
    end

    reg [7:0] out5611;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5611 = in0;
    end

    reg [7:0] out5612;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5612 = in0;
    end

    reg [7:0] out5613;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5613 = in0;
    end

    reg [7:0] out5614;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5614 = in0;
    end

    reg [7:0] out5615;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5615 = in0;
    end

    reg [7:0] out5616;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5616 = in0;
    end

    reg [7:0] out5617;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5617 = in0;
    end

    reg [7:0] out5618;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5618 = in0;
    end

    reg [7:0] out5619;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5619 = in0;
    end

    reg [7:0] out5620;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5620 = in0;
    end

    reg [7:0] out5621;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5621 = in0;
    end

    reg [7:0] out5622;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5622 = in0;
    end

    reg [7:0] out5623;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5623 = in0;
    end

    reg [7:0] out5624;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5624 = in0;
    end

    reg [7:0] out5625;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5625 = in0;
    end

    reg [7:0] out5626;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5626 = in0;
    end

    reg [7:0] out5627;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5627 = in0;
    end

    reg [7:0] out5628;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5628 = in0;
    end

    reg [7:0] out5629;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5629 = in0;
    end

    reg [7:0] out5630;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5630 = in0;
    end

    reg [7:0] out5631;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5631 = in0;
    end

    reg [7:0] out5632;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5632 = in0;
    end

    reg [7:0] out5633;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5633 = in0;
    end

    reg [7:0] out5634;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5634 = in0;
    end

    reg [7:0] out5635;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5635 = in0;
    end

    reg [7:0] out5636;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5636 = in0;
    end

    reg [7:0] out5637;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5637 = in0;
    end

    reg [7:0] out5638;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5638 = in0;
    end

    reg [7:0] out5639;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5639 = in0;
    end

    reg [7:0] out5640;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5640 = in0;
    end

    reg [7:0] out5641;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5641 = in0;
    end

    reg [7:0] out5642;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5642 = in0;
    end

    reg [7:0] out5643;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5643 = in0;
    end

    reg [7:0] out5644;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5644 = in0;
    end

    reg [7:0] out5645;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5645 = in0;
    end

    reg [7:0] out5646;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5646 = in0;
    end

    reg [7:0] out5647;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5647 = in0;
    end

    reg [7:0] out5648;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5648 = in0;
    end

    reg [7:0] out5649;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5649 = in0;
    end

    reg [7:0] out5650;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5650 = in0;
    end

    reg [7:0] out5651;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5651 = in0;
    end

    reg [7:0] out5652;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5652 = in0;
    end

    reg [7:0] out5653;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5653 = in0;
    end

    reg [7:0] out5654;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5654 = in0;
    end

    reg [7:0] out5655;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5655 = in0;
    end

    reg [7:0] out5656;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5656 = in0;
    end

    reg [7:0] out5657;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5657 = in0;
    end

    reg [7:0] out5658;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5658 = in0;
    end

    reg [7:0] out5659;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5659 = in0;
    end

    reg [7:0] out5660;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5660 = in0;
    end

    reg [7:0] out5661;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5661 = in0;
    end

    reg [7:0] out5662;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5662 = in0;
    end

    reg [7:0] out5663;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5663 = in0;
    end

    reg [7:0] out5664;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5664 = in0;
    end

    reg [7:0] out5665;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5665 = in0;
    end

    reg [7:0] out5666;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5666 = in0;
    end

    reg [7:0] out5667;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5667 = in0;
    end

    reg [7:0] out5668;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5668 = in0;
    end

    reg [7:0] out5669;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5669 = in0;
    end

    reg [7:0] out5670;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5670 = in0;
    end

    reg [7:0] out5671;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5671 = in0;
    end

    reg [7:0] out5672;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5672 = in0;
    end

    reg [7:0] out5673;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5673 = in0;
    end

    reg [7:0] out5674;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5674 = in0;
    end

    reg [7:0] out5675;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5675 = in0;
    end

    reg [7:0] out5676;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5676 = in0;
    end

    reg [7:0] out5677;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5677 = in0;
    end

    reg [7:0] out5678;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5678 = in0;
    end

    reg [7:0] out5679;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5679 = in0;
    end

    reg [7:0] out5680;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5680 = in0;
    end

    reg [7:0] out5681;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5681 = in0;
    end

    reg [7:0] out5682;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5682 = in0;
    end

    reg [7:0] out5683;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5683 = in0;
    end

    reg [7:0] out5684;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5684 = in0;
    end

    reg [7:0] out5685;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5685 = in0;
    end

    reg [7:0] out5686;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5686 = in0;
    end

    reg [7:0] out5687;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5687 = in0;
    end

    reg [7:0] out5688;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5688 = in0;
    end

    reg [7:0] out5689;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5689 = in0;
    end

    reg [7:0] out5690;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5690 = in0;
    end

    reg [7:0] out5691;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5691 = in0;
    end

    reg [7:0] out5692;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5692 = in0;
    end

    reg [7:0] out5693;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5693 = in0;
    end

    reg [7:0] out5694;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5694 = in0;
    end

    reg [7:0] out5695;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5695 = in0;
    end

    reg [7:0] out5696;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5696 = in0;
    end

    reg [7:0] out5697;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5697 = in0;
    end

    reg [7:0] out5698;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5698 = in0;
    end

    reg [7:0] out5699;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5699 = in0;
    end

    reg [7:0] out5700;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5700 = in0;
    end

    reg [7:0] out5701;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5701 = in0;
    end

    reg [7:0] out5702;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5702 = in0;
    end

    reg [7:0] out5703;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5703 = in0;
    end

    reg [7:0] out5704;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5704 = in0;
    end

    reg [7:0] out5705;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5705 = in0;
    end

    reg [7:0] out5706;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5706 = in0;
    end

    reg [7:0] out5707;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5707 = in0;
    end

    reg [7:0] out5708;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5708 = in0;
    end

    reg [7:0] out5709;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5709 = in0;
    end

    reg [7:0] out5710;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5710 = in0;
    end

    reg [7:0] out5711;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5711 = in0;
    end

    reg [7:0] out5712;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5712 = in0;
    end

    reg [7:0] out5713;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5713 = in0;
    end

    reg [7:0] out5714;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5714 = in0;
    end

    reg [7:0] out5715;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5715 = in0;
    end

    reg [7:0] out5716;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5716 = in0;
    end

    reg [7:0] out5717;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5717 = in0;
    end

    reg [7:0] out5718;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5718 = in0;
    end

    reg [7:0] out5719;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5719 = in0;
    end

    reg [7:0] out5720;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5720 = in0;
    end

    reg [7:0] out5721;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5721 = in0;
    end

    reg [7:0] out5722;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5722 = in0;
    end

    reg [7:0] out5723;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5723 = in0;
    end

    reg [7:0] out5724;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5724 = in0;
    end

    reg [7:0] out5725;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5725 = in0;
    end

    reg [7:0] out5726;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5726 = in0;
    end

    reg [7:0] out5727;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5727 = in0;
    end

    reg [7:0] out5728;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5728 = in0;
    end

    reg [7:0] out5729;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5729 = in0;
    end

    reg [7:0] out5730;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5730 = in0;
    end

    reg [7:0] out5731;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5731 = in0;
    end

    reg [7:0] out5732;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5732 = in0;
    end

    reg [7:0] out5733;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5733 = in0;
    end

    reg [7:0] out5734;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5734 = in0;
    end

    reg [7:0] out5735;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5735 = in0;
    end

    reg [7:0] out5736;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5736 = in0;
    end

    reg [7:0] out5737;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5737 = in0;
    end

    reg [7:0] out5738;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5738 = in0;
    end

    reg [7:0] out5739;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5739 = in0;
    end

    reg [7:0] out5740;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5740 = in0;
    end

    reg [7:0] out5741;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5741 = in0;
    end

    reg [7:0] out5742;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5742 = in0;
    end

    reg [7:0] out5743;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5743 = in0;
    end

    reg [7:0] out5744;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5744 = in0;
    end

    reg [7:0] out5745;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5745 = in0;
    end

    reg [7:0] out5746;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5746 = in0;
    end

    reg [7:0] out5747;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5747 = in0;
    end

    reg [7:0] out5748;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5748 = in0;
    end

    reg [7:0] out5749;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5749 = in0;
    end

    reg [7:0] out5750;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5750 = in0;
    end

    reg [7:0] out5751;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5751 = in0;
    end

    reg [7:0] out5752;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5752 = in0;
    end

    reg [7:0] out5753;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5753 = in0;
    end

    reg [7:0] out5754;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5754 = in0;
    end

    reg [7:0] out5755;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5755 = in0;
    end

    reg [7:0] out5756;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5756 = in0;
    end

    reg [7:0] out5757;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5757 = in0;
    end

    reg [7:0] out5758;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5758 = in0;
    end

    reg [7:0] out5759;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5759 = in0;
    end

    reg [7:0] out5760;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5760 = in0;
    end

    reg [7:0] out5761;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5761 = in0;
    end

    reg [7:0] out5762;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5762 = in0;
    end

    reg [7:0] out5763;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5763 = in0;
    end

    reg [7:0] out5764;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5764 = in0;
    end

    reg [7:0] out5765;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5765 = in0;
    end

    reg [7:0] out5766;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5766 = in0;
    end

    reg [7:0] out5767;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5767 = in0;
    end

    reg [7:0] out5768;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5768 = in0;
    end

    reg [7:0] out5769;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5769 = in0;
    end

    reg [7:0] out5770;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5770 = in0;
    end

    reg [7:0] out5771;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5771 = in0;
    end

    reg [7:0] out5772;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5772 = in0;
    end

    reg [7:0] out5773;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5773 = in0;
    end

    reg [7:0] out5774;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5774 = in0;
    end

    reg [7:0] out5775;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5775 = in0;
    end

    reg [7:0] out5776;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5776 = in0;
    end

    reg [7:0] out5777;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5777 = in0;
    end

    reg [7:0] out5778;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5778 = in0;
    end

    reg [7:0] out5779;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5779 = in0;
    end

    reg [7:0] out5780;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5780 = in0;
    end

    reg [7:0] out5781;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5781 = in0;
    end

    reg [7:0] out5782;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5782 = in0;
    end

    reg [7:0] out5783;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5783 = in0;
    end

    reg [7:0] out5784;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5784 = in0;
    end

    reg [7:0] out5785;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5785 = in0;
    end

    reg [7:0] out5786;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5786 = in0;
    end

    reg [7:0] out5787;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5787 = in0;
    end

    reg [7:0] out5788;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5788 = in0;
    end

    reg [7:0] out5789;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5789 = in0;
    end

    reg [7:0] out5790;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5790 = in0;
    end

    reg [7:0] out5791;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5791 = in0;
    end

    reg [7:0] out5792;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5792 = in0;
    end

    reg [7:0] out5793;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5793 = in0;
    end

    reg [7:0] out5794;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5794 = in0;
    end

    reg [7:0] out5795;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5795 = in0;
    end

    reg [7:0] out5796;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5796 = in0;
    end

    reg [7:0] out5797;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5797 = in0;
    end

    reg [7:0] out5798;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5798 = in0;
    end

    reg [7:0] out5799;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5799 = in0;
    end

    reg [7:0] out5800;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5800 = in0;
    end

    reg [7:0] out5801;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5801 = in0;
    end

    reg [7:0] out5802;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5802 = in0;
    end

    reg [7:0] out5803;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5803 = in0;
    end

    reg [7:0] out5804;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5804 = in0;
    end

    reg [7:0] out5805;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5805 = in0;
    end

    reg [7:0] out5806;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5806 = in0;
    end

    reg [7:0] out5807;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5807 = in0;
    end

    reg [7:0] out5808;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5808 = in0;
    end

    reg [7:0] out5809;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5809 = in0;
    end

    reg [7:0] out5810;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5810 = in0;
    end

    reg [7:0] out5811;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5811 = in0;
    end

    reg [7:0] out5812;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5812 = in0;
    end

    reg [7:0] out5813;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5813 = in0;
    end

    reg [7:0] out5814;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5814 = in0;
    end

    reg [7:0] out5815;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5815 = in0;
    end

    reg [7:0] out5816;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5816 = in0;
    end

    reg [7:0] out5817;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5817 = in0;
    end

    reg [7:0] out5818;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5818 = in0;
    end

    reg [7:0] out5819;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5819 = in0;
    end

    reg [7:0] out5820;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5820 = in0;
    end

    reg [7:0] out5821;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5821 = in0;
    end

    reg [7:0] out5822;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5822 = in0;
    end

    reg [7:0] out5823;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5823 = in0;
    end

    reg [7:0] out5824;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5824 = in0;
    end

    reg [7:0] out5825;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5825 = in0;
    end

    reg [7:0] out5826;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5826 = in0;
    end

    reg [7:0] out5827;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5827 = in0;
    end

    reg [7:0] out5828;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5828 = in0;
    end

    reg [7:0] out5829;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5829 = in0;
    end

    reg [7:0] out5830;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5830 = in0;
    end

    reg [7:0] out5831;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5831 = in0;
    end

    reg [7:0] out5832;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5832 = in0;
    end

    reg [7:0] out5833;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5833 = in0;
    end

    reg [7:0] out5834;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5834 = in0;
    end

    reg [7:0] out5835;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5835 = in0;
    end

    reg [7:0] out5836;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5836 = in0;
    end

    reg [7:0] out5837;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5837 = in0;
    end

    reg [7:0] out5838;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5838 = in0;
    end

    reg [7:0] out5839;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5839 = in0;
    end

    reg [7:0] out5840;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5840 = in0;
    end

    reg [7:0] out5841;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5841 = in0;
    end

    reg [7:0] out5842;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5842 = in0;
    end

    reg [7:0] out5843;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5843 = in0;
    end

    reg [7:0] out5844;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5844 = in0;
    end

    reg [7:0] out5845;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5845 = in0;
    end

    reg [7:0] out5846;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5846 = in0;
    end

    reg [7:0] out5847;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5847 = in0;
    end

    reg [7:0] out5848;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5848 = in0;
    end

    reg [7:0] out5849;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5849 = in0;
    end

    reg [7:0] out5850;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5850 = in0;
    end

    reg [7:0] out5851;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5851 = in0;
    end

    reg [7:0] out5852;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5852 = in0;
    end

    reg [7:0] out5853;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5853 = in0;
    end

    reg [7:0] out5854;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5854 = in0;
    end

    reg [7:0] out5855;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5855 = in0;
    end

    reg [7:0] out5856;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5856 = in0;
    end

    reg [7:0] out5857;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5857 = in0;
    end

    reg [7:0] out5858;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5858 = in0;
    end

    reg [7:0] out5859;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5859 = in0;
    end

    reg [7:0] out5860;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5860 = in0;
    end

    reg [7:0] out5861;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5861 = in0;
    end

    reg [7:0] out5862;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5862 = in0;
    end

    reg [7:0] out5863;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5863 = in0;
    end

    reg [7:0] out5864;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5864 = in0;
    end

    reg [7:0] out5865;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5865 = in0;
    end

    reg [7:0] out5866;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5866 = in0;
    end

    reg [7:0] out5867;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5867 = in0;
    end

    reg [7:0] out5868;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5868 = in0;
    end

    reg [7:0] out5869;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5869 = in0;
    end

    reg [7:0] out5870;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5870 = in0;
    end

    reg [7:0] out5871;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5871 = in0;
    end

    reg [7:0] out5872;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5872 = in0;
    end

    reg [7:0] out5873;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5873 = in0;
    end

    reg [7:0] out5874;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5874 = in0;
    end

    reg [7:0] out5875;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5875 = in0;
    end

    reg [7:0] out5876;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5876 = in0;
    end

    reg [7:0] out5877;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5877 = in0;
    end

    reg [7:0] out5878;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5878 = in0;
    end

    reg [7:0] out5879;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5879 = in0;
    end

    reg [7:0] out5880;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5880 = in0;
    end

    reg [7:0] out5881;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5881 = in0;
    end

    reg [7:0] out5882;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5882 = in0;
    end

    reg [7:0] out5883;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5883 = in0;
    end

    reg [7:0] out5884;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5884 = in0;
    end

    reg [7:0] out5885;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5885 = in0;
    end

    reg [7:0] out5886;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5886 = in0;
    end

    reg [7:0] out5887;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5887 = in0;
    end

    reg [7:0] out5888;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5888 = in0;
    end

    reg [7:0] out5889;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5889 = in0;
    end

    reg [7:0] out5890;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5890 = in0;
    end

    reg [7:0] out5891;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5891 = in0;
    end

    reg [7:0] out5892;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5892 = in0;
    end

    reg [7:0] out5893;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5893 = in0;
    end

    reg [7:0] out5894;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5894 = in0;
    end

    reg [7:0] out5895;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5895 = in0;
    end

    reg [7:0] out5896;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5896 = in0;
    end

    reg [7:0] out5897;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5897 = in0;
    end

    reg [7:0] out5898;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5898 = in0;
    end

    reg [7:0] out5899;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5899 = in0;
    end

    reg [7:0] out5900;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5900 = in0;
    end

    reg [7:0] out5901;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5901 = in0;
    end

    reg [7:0] out5902;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5902 = in0;
    end

    reg [7:0] out5903;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5903 = in0;
    end

    reg [7:0] out5904;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5904 = in0;
    end

    reg [7:0] out5905;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5905 = in0;
    end

    reg [7:0] out5906;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5906 = in0;
    end

    reg [7:0] out5907;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5907 = in0;
    end

    reg [7:0] out5908;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5908 = in0;
    end

    reg [7:0] out5909;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5909 = in0;
    end

    reg [7:0] out5910;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5910 = in0;
    end

    reg [7:0] out5911;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5911 = in0;
    end

    reg [7:0] out5912;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5912 = in0;
    end

    reg [7:0] out5913;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5913 = in0;
    end

    reg [7:0] out5914;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5914 = in0;
    end

    reg [7:0] out5915;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5915 = in0;
    end

    reg [7:0] out5916;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5916 = in0;
    end

    reg [7:0] out5917;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5917 = in0;
    end

    reg [7:0] out5918;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5918 = in0;
    end

    reg [7:0] out5919;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5919 = in0;
    end

    reg [7:0] out5920;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5920 = in0;
    end

    reg [7:0] out5921;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5921 = in0;
    end

    reg [7:0] out5922;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5922 = in0;
    end

    reg [7:0] out5923;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5923 = in0;
    end

    reg [7:0] out5924;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5924 = in0;
    end

    reg [7:0] out5925;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5925 = in0;
    end

    reg [7:0] out5926;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5926 = in0;
    end

    reg [7:0] out5927;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5927 = in0;
    end

    reg [7:0] out5928;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5928 = in0;
    end

    reg [7:0] out5929;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5929 = in0;
    end

    reg [7:0] out5930;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5930 = in0;
    end

    reg [7:0] out5931;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5931 = in0;
    end

    reg [7:0] out5932;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5932 = in0;
    end

    reg [7:0] out5933;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5933 = in0;
    end

    reg [7:0] out5934;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5934 = in0;
    end

    reg [7:0] out5935;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5935 = in0;
    end

    reg [7:0] out5936;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5936 = in0;
    end

    reg [7:0] out5937;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5937 = in0;
    end

    reg [7:0] out5938;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5938 = in0;
    end

    reg [7:0] out5939;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5939 = in0;
    end

    reg [7:0] out5940;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5940 = in0;
    end

    reg [7:0] out5941;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5941 = in0;
    end

    reg [7:0] out5942;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5942 = in0;
    end

    reg [7:0] out5943;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5943 = in0;
    end

    reg [7:0] out5944;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5944 = in0;
    end

    reg [7:0] out5945;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5945 = in0;
    end

    reg [7:0] out5946;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5946 = in0;
    end

    reg [7:0] out5947;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5947 = in0;
    end

    reg [7:0] out5948;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5948 = in0;
    end

    reg [7:0] out5949;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5949 = in0;
    end

    reg [7:0] out5950;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5950 = in0;
    end

    reg [7:0] out5951;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5951 = in0;
    end

    reg [7:0] out5952;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5952 = in0;
    end

    reg [7:0] out5953;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5953 = in0;
    end

    reg [7:0] out5954;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5954 = in0;
    end

    reg [7:0] out5955;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5955 = in0;
    end

    reg [7:0] out5956;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5956 = in0;
    end

    reg [7:0] out5957;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5957 = in0;
    end

    reg [7:0] out5958;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5958 = in0;
    end

    reg [7:0] out5959;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5959 = in0;
    end

    reg [7:0] out5960;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5960 = in0;
    end

    reg [7:0] out5961;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5961 = in0;
    end

    reg [7:0] out5962;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5962 = in0;
    end

    reg [7:0] out5963;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5963 = in0;
    end

    reg [7:0] out5964;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5964 = in0;
    end

    reg [7:0] out5965;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5965 = in0;
    end

    reg [7:0] out5966;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5966 = in0;
    end

    reg [7:0] out5967;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5967 = in0;
    end

    reg [7:0] out5968;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5968 = in0;
    end

    reg [7:0] out5969;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5969 = in0;
    end

    reg [7:0] out5970;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5970 = in0;
    end

    reg [7:0] out5971;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5971 = in0;
    end

    reg [7:0] out5972;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5972 = in0;
    end

    reg [7:0] out5973;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5973 = in0;
    end

    reg [7:0] out5974;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5974 = in0;
    end

    reg [7:0] out5975;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5975 = in0;
    end

    reg [7:0] out5976;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5976 = in0;
    end

    reg [7:0] out5977;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5977 = in0;
    end

    reg [7:0] out5978;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5978 = in0;
    end

    reg [7:0] out5979;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5979 = in0;
    end

    reg [7:0] out5980;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5980 = in0;
    end

    reg [7:0] out5981;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5981 = in0;
    end

    reg [7:0] out5982;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5982 = in0;
    end

    reg [7:0] out5983;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5983 = in0;
    end

    reg [7:0] out5984;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5984 = in0;
    end

    reg [7:0] out5985;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5985 = in0;
    end

    reg [7:0] out5986;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5986 = in0;
    end

    reg [7:0] out5987;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5987 = in0;
    end

    reg [7:0] out5988;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5988 = in0;
    end

    reg [7:0] out5989;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5989 = in0;
    end

    reg [7:0] out5990;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5990 = in0;
    end

    reg [7:0] out5991;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5991 = in0;
    end

    reg [7:0] out5992;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5992 = in0;
    end

    reg [7:0] out5993;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5993 = in0;
    end

    reg [7:0] out5994;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5994 = in0;
    end

    reg [7:0] out5995;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5995 = in0;
    end

    reg [7:0] out5996;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5996 = in0;
    end

    reg [7:0] out5997;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5997 = in0;
    end

    reg [7:0] out5998;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5998 = in0;
    end

    reg [7:0] out5999;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out5999 = in0;
    end

    reg [7:0] out6000;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6000 = in0;
    end

    reg [7:0] out6001;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6001 = in0;
    end

    reg [7:0] out6002;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6002 = in0;
    end

    reg [7:0] out6003;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6003 = in0;
    end

    reg [7:0] out6004;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6004 = in0;
    end

    reg [7:0] out6005;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6005 = in0;
    end

    reg [7:0] out6006;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6006 = in0;
    end

    reg [7:0] out6007;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6007 = in0;
    end

    reg [7:0] out6008;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6008 = in0;
    end

    reg [7:0] out6009;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6009 = in0;
    end

    reg [7:0] out6010;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6010 = in0;
    end

    reg [7:0] out6011;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6011 = in0;
    end

    reg [7:0] out6012;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6012 = in0;
    end

    reg [7:0] out6013;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6013 = in0;
    end

    reg [7:0] out6014;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6014 = in0;
    end

    reg [7:0] out6015;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6015 = in0;
    end

    reg [7:0] out6016;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6016 = in0;
    end

    reg [7:0] out6017;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6017 = in0;
    end

    reg [7:0] out6018;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6018 = in0;
    end

    reg [7:0] out6019;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6019 = in0;
    end

    reg [7:0] out6020;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6020 = in0;
    end

    reg [7:0] out6021;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6021 = in0;
    end

    reg [7:0] out6022;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6022 = in0;
    end

    reg [7:0] out6023;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6023 = in0;
    end

    reg [7:0] out6024;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6024 = in0;
    end

    reg [7:0] out6025;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6025 = in0;
    end

    reg [7:0] out6026;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6026 = in0;
    end

    reg [7:0] out6027;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6027 = in0;
    end

    reg [7:0] out6028;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6028 = in0;
    end

    reg [7:0] out6029;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6029 = in0;
    end

    reg [7:0] out6030;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6030 = in0;
    end

    reg [7:0] out6031;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6031 = in0;
    end

    reg [7:0] out6032;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6032 = in0;
    end

    reg [7:0] out6033;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6033 = in0;
    end

    reg [7:0] out6034;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6034 = in0;
    end

    reg [7:0] out6035;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6035 = in0;
    end

    reg [7:0] out6036;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6036 = in0;
    end

    reg [7:0] out6037;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6037 = in0;
    end

    reg [7:0] out6038;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6038 = in0;
    end

    reg [7:0] out6039;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6039 = in0;
    end

    reg [7:0] out6040;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6040 = in0;
    end

    reg [7:0] out6041;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6041 = in0;
    end

    reg [7:0] out6042;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6042 = in0;
    end

    reg [7:0] out6043;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6043 = in0;
    end

    reg [7:0] out6044;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6044 = in0;
    end

    reg [7:0] out6045;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6045 = in0;
    end

    reg [7:0] out6046;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6046 = in0;
    end

    reg [7:0] out6047;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6047 = in0;
    end

    reg [7:0] out6048;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6048 = in0;
    end

    reg [7:0] out6049;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6049 = in0;
    end

    reg [7:0] out6050;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6050 = in0;
    end

    reg [7:0] out6051;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6051 = in0;
    end

    reg [7:0] out6052;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6052 = in0;
    end

    reg [7:0] out6053;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6053 = in0;
    end

    reg [7:0] out6054;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6054 = in0;
    end

    reg [7:0] out6055;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6055 = in0;
    end

    reg [7:0] out6056;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6056 = in0;
    end

    reg [7:0] out6057;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6057 = in0;
    end

    reg [7:0] out6058;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6058 = in0;
    end

    reg [7:0] out6059;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6059 = in0;
    end

    reg [7:0] out6060;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6060 = in0;
    end

    reg [7:0] out6061;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6061 = in0;
    end

    reg [7:0] out6062;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6062 = in0;
    end

    reg [7:0] out6063;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6063 = in0;
    end

    reg [7:0] out6064;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6064 = in0;
    end

    reg [7:0] out6065;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6065 = in0;
    end

    reg [7:0] out6066;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6066 = in0;
    end

    reg [7:0] out6067;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6067 = in0;
    end

    reg [7:0] out6068;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6068 = in0;
    end

    reg [7:0] out6069;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6069 = in0;
    end

    reg [7:0] out6070;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6070 = in0;
    end

    reg [7:0] out6071;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6071 = in0;
    end

    reg [7:0] out6072;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6072 = in0;
    end

    reg [7:0] out6073;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6073 = in0;
    end

    reg [7:0] out6074;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6074 = in0;
    end

    reg [7:0] out6075;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6075 = in0;
    end

    reg [7:0] out6076;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6076 = in0;
    end

    reg [7:0] out6077;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6077 = in0;
    end

    reg [7:0] out6078;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6078 = in0;
    end

    reg [7:0] out6079;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6079 = in0;
    end

    reg [7:0] out6080;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6080 = in0;
    end

    reg [7:0] out6081;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6081 = in0;
    end

    reg [7:0] out6082;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6082 = in0;
    end

    reg [7:0] out6083;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6083 = in0;
    end

    reg [7:0] out6084;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6084 = in0;
    end

    reg [7:0] out6085;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6085 = in0;
    end

    reg [7:0] out6086;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6086 = in0;
    end

    reg [7:0] out6087;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6087 = in0;
    end

    reg [7:0] out6088;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6088 = in0;
    end

    reg [7:0] out6089;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6089 = in0;
    end

    reg [7:0] out6090;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6090 = in0;
    end

    reg [7:0] out6091;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6091 = in0;
    end

    reg [7:0] out6092;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6092 = in0;
    end

    reg [7:0] out6093;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6093 = in0;
    end

    reg [7:0] out6094;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6094 = in0;
    end

    reg [7:0] out6095;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6095 = in0;
    end

    reg [7:0] out6096;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6096 = in0;
    end

    reg [7:0] out6097;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6097 = in0;
    end

    reg [7:0] out6098;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6098 = in0;
    end

    reg [7:0] out6099;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6099 = in0;
    end

    reg [7:0] out6100;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6100 = in0;
    end

    reg [7:0] out6101;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6101 = in0;
    end

    reg [7:0] out6102;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6102 = in0;
    end

    reg [7:0] out6103;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6103 = in0;
    end

    reg [7:0] out6104;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6104 = in0;
    end

    reg [7:0] out6105;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6105 = in0;
    end

    reg [7:0] out6106;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6106 = in0;
    end

    reg [7:0] out6107;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6107 = in0;
    end

    reg [7:0] out6108;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6108 = in0;
    end

    reg [7:0] out6109;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6109 = in0;
    end

    reg [7:0] out6110;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6110 = in0;
    end

    reg [7:0] out6111;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6111 = in0;
    end

    reg [7:0] out6112;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6112 = in0;
    end

    reg [7:0] out6113;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6113 = in0;
    end

    reg [7:0] out6114;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6114 = in0;
    end

    reg [7:0] out6115;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6115 = in0;
    end

    reg [7:0] out6116;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6116 = in0;
    end

    reg [7:0] out6117;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6117 = in0;
    end

    reg [7:0] out6118;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6118 = in0;
    end

    reg [7:0] out6119;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6119 = in0;
    end

    reg [7:0] out6120;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6120 = in0;
    end

    reg [7:0] out6121;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6121 = in0;
    end

    reg [7:0] out6122;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6122 = in0;
    end

    reg [7:0] out6123;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6123 = in0;
    end

    reg [7:0] out6124;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6124 = in0;
    end

    reg [7:0] out6125;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6125 = in0;
    end

    reg [7:0] out6126;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6126 = in0;
    end

    reg [7:0] out6127;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6127 = in0;
    end

    reg [7:0] out6128;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6128 = in0;
    end

    reg [7:0] out6129;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6129 = in0;
    end

    reg [7:0] out6130;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6130 = in0;
    end

    reg [7:0] out6131;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6131 = in0;
    end

    reg [7:0] out6132;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6132 = in0;
    end

    reg [7:0] out6133;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6133 = in0;
    end

    reg [7:0] out6134;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6134 = in0;
    end

    reg [7:0] out6135;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6135 = in0;
    end

    reg [7:0] out6136;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6136 = in0;
    end

    reg [7:0] out6137;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6137 = in0;
    end

    reg [7:0] out6138;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6138 = in0;
    end

    reg [7:0] out6139;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6139 = in0;
    end

    reg [7:0] out6140;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6140 = in0;
    end

    reg [7:0] out6141;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6141 = in0;
    end

    reg [7:0] out6142;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6142 = in0;
    end

    reg [7:0] out6143;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6143 = in0;
    end

    reg [7:0] out6144;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6144 = in0;
    end

    reg [7:0] out6145;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6145 = in0;
    end

    reg [7:0] out6146;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6146 = in0;
    end

    reg [7:0] out6147;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6147 = in0;
    end

    reg [7:0] out6148;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6148 = in0;
    end

    reg [7:0] out6149;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6149 = in0;
    end

    reg [7:0] out6150;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6150 = in0;
    end

    reg [7:0] out6151;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6151 = in0;
    end

    reg [7:0] out6152;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6152 = in0;
    end

    reg [7:0] out6153;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6153 = in0;
    end

    reg [7:0] out6154;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6154 = in0;
    end

    reg [7:0] out6155;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6155 = in0;
    end

    reg [7:0] out6156;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6156 = in0;
    end

    reg [7:0] out6157;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6157 = in0;
    end

    reg [7:0] out6158;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6158 = in0;
    end

    reg [7:0] out6159;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6159 = in0;
    end

    reg [7:0] out6160;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6160 = in0;
    end

    reg [7:0] out6161;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6161 = in0;
    end

    reg [7:0] out6162;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6162 = in0;
    end

    reg [7:0] out6163;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6163 = in0;
    end

    reg [7:0] out6164;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6164 = in0;
    end

    reg [7:0] out6165;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6165 = in0;
    end

    reg [7:0] out6166;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6166 = in0;
    end

    reg [7:0] out6167;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6167 = in0;
    end

    reg [7:0] out6168;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6168 = in0;
    end

    reg [7:0] out6169;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6169 = in0;
    end

    reg [7:0] out6170;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6170 = in0;
    end

    reg [7:0] out6171;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6171 = in0;
    end

    reg [7:0] out6172;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6172 = in0;
    end

    reg [7:0] out6173;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6173 = in0;
    end

    reg [7:0] out6174;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6174 = in0;
    end

    reg [7:0] out6175;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6175 = in0;
    end

    reg [7:0] out6176;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6176 = in0;
    end

    reg [7:0] out6177;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6177 = in0;
    end

    reg [7:0] out6178;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6178 = in0;
    end

    reg [7:0] out6179;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6179 = in0;
    end

    reg [7:0] out6180;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6180 = in0;
    end

    reg [7:0] out6181;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6181 = in0;
    end

    reg [7:0] out6182;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6182 = in0;
    end

    reg [7:0] out6183;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6183 = in0;
    end

    reg [7:0] out6184;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6184 = in0;
    end

    reg [7:0] out6185;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6185 = in0;
    end

    reg [7:0] out6186;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6186 = in0;
    end

    reg [7:0] out6187;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6187 = in0;
    end

    reg [7:0] out6188;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6188 = in0;
    end

    reg [7:0] out6189;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6189 = in0;
    end

    reg [7:0] out6190;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6190 = in0;
    end

    reg [7:0] out6191;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6191 = in0;
    end

    reg [7:0] out6192;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6192 = in0;
    end

    reg [7:0] out6193;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6193 = in0;
    end

    reg [7:0] out6194;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6194 = in0;
    end

    reg [7:0] out6195;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6195 = in0;
    end

    reg [7:0] out6196;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6196 = in0;
    end

    reg [7:0] out6197;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6197 = in0;
    end

    reg [7:0] out6198;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6198 = in0;
    end

    reg [7:0] out6199;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6199 = in0;
    end

    reg [7:0] out6200;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6200 = in0;
    end

    reg [7:0] out6201;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6201 = in0;
    end

    reg [7:0] out6202;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6202 = in0;
    end

    reg [7:0] out6203;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6203 = in0;
    end

    reg [7:0] out6204;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6204 = in0;
    end

    reg [7:0] out6205;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6205 = in0;
    end

    reg [7:0] out6206;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6206 = in0;
    end

    reg [7:0] out6207;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6207 = in0;
    end

    reg [7:0] out6208;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6208 = in0;
    end

    reg [7:0] out6209;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6209 = in0;
    end

    reg [7:0] out6210;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6210 = in0;
    end

    reg [7:0] out6211;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6211 = in0;
    end

    reg [7:0] out6212;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6212 = in0;
    end

    reg [7:0] out6213;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6213 = in0;
    end

    reg [7:0] out6214;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6214 = in0;
    end

    reg [7:0] out6215;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6215 = in0;
    end

    reg [7:0] out6216;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6216 = in0;
    end

    reg [7:0] out6217;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6217 = in0;
    end

    reg [7:0] out6218;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6218 = in0;
    end

    reg [7:0] out6219;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6219 = in0;
    end

    reg [7:0] out6220;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6220 = in0;
    end

    reg [7:0] out6221;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6221 = in0;
    end

    reg [7:0] out6222;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6222 = in0;
    end

    reg [7:0] out6223;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6223 = in0;
    end

    reg [7:0] out6224;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6224 = in0;
    end

    reg [7:0] out6225;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6225 = in0;
    end

    reg [7:0] out6226;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6226 = in0;
    end

    reg [7:0] out6227;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6227 = in0;
    end

    reg [7:0] out6228;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6228 = in0;
    end

    reg [7:0] out6229;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6229 = in0;
    end

    reg [7:0] out6230;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6230 = in0;
    end

    reg [7:0] out6231;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6231 = in0;
    end

    reg [7:0] out6232;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6232 = in0;
    end

    reg [7:0] out6233;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6233 = in0;
    end

    reg [7:0] out6234;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6234 = in0;
    end

    reg [7:0] out6235;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6235 = in0;
    end

    reg [7:0] out6236;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6236 = in0;
    end

    reg [7:0] out6237;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6237 = in0;
    end

    reg [7:0] out6238;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6238 = in0;
    end

    reg [7:0] out6239;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6239 = in0;
    end

    reg [7:0] out6240;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6240 = in0;
    end

    reg [7:0] out6241;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6241 = in0;
    end

    reg [7:0] out6242;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6242 = in0;
    end

    reg [7:0] out6243;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6243 = in0;
    end

    reg [7:0] out6244;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6244 = in0;
    end

    reg [7:0] out6245;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6245 = in0;
    end

    reg [7:0] out6246;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6246 = in0;
    end

    reg [7:0] out6247;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6247 = in0;
    end

    reg [7:0] out6248;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6248 = in0;
    end

    reg [7:0] out6249;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6249 = in0;
    end

    reg [7:0] out6250;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6250 = in0;
    end

    reg [7:0] out6251;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6251 = in0;
    end

    reg [7:0] out6252;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6252 = in0;
    end

    reg [7:0] out6253;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6253 = in0;
    end

    reg [7:0] out6254;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6254 = in0;
    end

    reg [7:0] out6255;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6255 = in0;
    end

    reg [7:0] out6256;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6256 = in0;
    end

    reg [7:0] out6257;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6257 = in0;
    end

    reg [7:0] out6258;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6258 = in0;
    end

    reg [7:0] out6259;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6259 = in0;
    end

    reg [7:0] out6260;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6260 = in0;
    end

    reg [7:0] out6261;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6261 = in0;
    end

    reg [7:0] out6262;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6262 = in0;
    end

    reg [7:0] out6263;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6263 = in0;
    end

    reg [7:0] out6264;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6264 = in0;
    end

    reg [7:0] out6265;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6265 = in0;
    end

    reg [7:0] out6266;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6266 = in0;
    end

    reg [7:0] out6267;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6267 = in0;
    end

    reg [7:0] out6268;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6268 = in0;
    end

    reg [7:0] out6269;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6269 = in0;
    end

    reg [7:0] out6270;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6270 = in0;
    end

    reg [7:0] out6271;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6271 = in0;
    end

    reg [7:0] out6272;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6272 = in0;
    end

    reg [7:0] out6273;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6273 = in0;
    end

    reg [7:0] out6274;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6274 = in0;
    end

    reg [7:0] out6275;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6275 = in0;
    end

    reg [7:0] out6276;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6276 = in0;
    end

    reg [7:0] out6277;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6277 = in0;
    end

    reg [7:0] out6278;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6278 = in0;
    end

    reg [7:0] out6279;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6279 = in0;
    end

    reg [7:0] out6280;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6280 = in0;
    end

    reg [7:0] out6281;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6281 = in0;
    end

    reg [7:0] out6282;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6282 = in0;
    end

    reg [7:0] out6283;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6283 = in0;
    end

    reg [7:0] out6284;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6284 = in0;
    end

    reg [7:0] out6285;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6285 = in0;
    end

    reg [7:0] out6286;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6286 = in0;
    end

    reg [7:0] out6287;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6287 = in0;
    end

    reg [7:0] out6288;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6288 = in0;
    end

    reg [7:0] out6289;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6289 = in0;
    end

    reg [7:0] out6290;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6290 = in0;
    end

    reg [7:0] out6291;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6291 = in0;
    end

    reg [7:0] out6292;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6292 = in0;
    end

    reg [7:0] out6293;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6293 = in0;
    end

    reg [7:0] out6294;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6294 = in0;
    end

    reg [7:0] out6295;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6295 = in0;
    end

    reg [7:0] out6296;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6296 = in0;
    end

    reg [7:0] out6297;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6297 = in0;
    end

    reg [7:0] out6298;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6298 = in0;
    end

    reg [7:0] out6299;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6299 = in0;
    end

    reg [7:0] out6300;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6300 = in0;
    end

    reg [7:0] out6301;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6301 = in0;
    end

    reg [7:0] out6302;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6302 = in0;
    end

    reg [7:0] out6303;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6303 = in0;
    end

    reg [7:0] out6304;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6304 = in0;
    end

    reg [7:0] out6305;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6305 = in0;
    end

    reg [7:0] out6306;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6306 = in0;
    end

    reg [7:0] out6307;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6307 = in0;
    end

    reg [7:0] out6308;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6308 = in0;
    end

    reg [7:0] out6309;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6309 = in0;
    end

    reg [7:0] out6310;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6310 = in0;
    end

    reg [7:0] out6311;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6311 = in0;
    end

    reg [7:0] out6312;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6312 = in0;
    end

    reg [7:0] out6313;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6313 = in0;
    end

    reg [7:0] out6314;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6314 = in0;
    end

    reg [7:0] out6315;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6315 = in0;
    end

    reg [7:0] out6316;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6316 = in0;
    end

    reg [7:0] out6317;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6317 = in0;
    end

    reg [7:0] out6318;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6318 = in0;
    end

    reg [7:0] out6319;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6319 = in0;
    end

    reg [7:0] out6320;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6320 = in0;
    end

    reg [7:0] out6321;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6321 = in0;
    end

    reg [7:0] out6322;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6322 = in0;
    end

    reg [7:0] out6323;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6323 = in0;
    end

    reg [7:0] out6324;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6324 = in0;
    end

    reg [7:0] out6325;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6325 = in0;
    end

    reg [7:0] out6326;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6326 = in0;
    end

    reg [7:0] out6327;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6327 = in0;
    end

    reg [7:0] out6328;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6328 = in0;
    end

    reg [7:0] out6329;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6329 = in0;
    end

    reg [7:0] out6330;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6330 = in0;
    end

    reg [7:0] out6331;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6331 = in0;
    end

    reg [7:0] out6332;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6332 = in0;
    end

    reg [7:0] out6333;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6333 = in0;
    end

    reg [7:0] out6334;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6334 = in0;
    end

    reg [7:0] out6335;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6335 = in0;
    end

    reg [7:0] out6336;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6336 = in0;
    end

    reg [7:0] out6337;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6337 = in0;
    end

    reg [7:0] out6338;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6338 = in0;
    end

    reg [7:0] out6339;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6339 = in0;
    end

    reg [7:0] out6340;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6340 = in0;
    end

    reg [7:0] out6341;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6341 = in0;
    end

    reg [7:0] out6342;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6342 = in0;
    end

    reg [7:0] out6343;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6343 = in0;
    end

    reg [7:0] out6344;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6344 = in0;
    end

    reg [7:0] out6345;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6345 = in0;
    end

    reg [7:0] out6346;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6346 = in0;
    end

    reg [7:0] out6347;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6347 = in0;
    end

    reg [7:0] out6348;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6348 = in0;
    end

    reg [7:0] out6349;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6349 = in0;
    end

    reg [7:0] out6350;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6350 = in0;
    end

    reg [7:0] out6351;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6351 = in0;
    end

    reg [7:0] out6352;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6352 = in0;
    end

    reg [7:0] out6353;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6353 = in0;
    end

    reg [7:0] out6354;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6354 = in0;
    end

    reg [7:0] out6355;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6355 = in0;
    end

    reg [7:0] out6356;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6356 = in0;
    end

    reg [7:0] out6357;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6357 = in0;
    end

    reg [7:0] out6358;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6358 = in0;
    end

    reg [7:0] out6359;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6359 = in0;
    end

    reg [7:0] out6360;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6360 = in0;
    end

    reg [7:0] out6361;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6361 = in0;
    end

    reg [7:0] out6362;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6362 = in0;
    end

    reg [7:0] out6363;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6363 = in0;
    end

    reg [7:0] out6364;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6364 = in0;
    end

    reg [7:0] out6365;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6365 = in0;
    end

    reg [7:0] out6366;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6366 = in0;
    end

    reg [7:0] out6367;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6367 = in0;
    end

    reg [7:0] out6368;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6368 = in0;
    end

    reg [7:0] out6369;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6369 = in0;
    end

    reg [7:0] out6370;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6370 = in0;
    end

    reg [7:0] out6371;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6371 = in0;
    end

    reg [7:0] out6372;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6372 = in0;
    end

    reg [7:0] out6373;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6373 = in0;
    end

    reg [7:0] out6374;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6374 = in0;
    end

    reg [7:0] out6375;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6375 = in0;
    end

    reg [7:0] out6376;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6376 = in0;
    end

    reg [7:0] out6377;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6377 = in0;
    end

    reg [7:0] out6378;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6378 = in0;
    end

    reg [7:0] out6379;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6379 = in0;
    end

    reg [7:0] out6380;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6380 = in0;
    end

    reg [7:0] out6381;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6381 = in0;
    end

    reg [7:0] out6382;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6382 = in0;
    end

    reg [7:0] out6383;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6383 = in0;
    end

    reg [7:0] out6384;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6384 = in0;
    end

    reg [7:0] out6385;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6385 = in0;
    end

    reg [7:0] out6386;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6386 = in0;
    end

    reg [7:0] out6387;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6387 = in0;
    end

    reg [7:0] out6388;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6388 = in0;
    end

    reg [7:0] out6389;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6389 = in0;
    end

    reg [7:0] out6390;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6390 = in0;
    end

    reg [7:0] out6391;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6391 = in0;
    end

    reg [7:0] out6392;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6392 = in0;
    end

    reg [7:0] out6393;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6393 = in0;
    end

    reg [7:0] out6394;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6394 = in0;
    end

    reg [7:0] out6395;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6395 = in0;
    end

    reg [7:0] out6396;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6396 = in0;
    end

    reg [7:0] out6397;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6397 = in0;
    end

    reg [7:0] out6398;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6398 = in0;
    end

    reg [7:0] out6399;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6399 = in0;
    end

    reg [7:0] out6400;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6400 = in0;
    end

    reg [7:0] out6401;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6401 = in0;
    end

    reg [7:0] out6402;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6402 = in0;
    end

    reg [7:0] out6403;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6403 = in0;
    end

    reg [7:0] out6404;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6404 = in0;
    end

    reg [7:0] out6405;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6405 = in0;
    end

    reg [7:0] out6406;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6406 = in0;
    end

    reg [7:0] out6407;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6407 = in0;
    end

    reg [7:0] out6408;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6408 = in0;
    end

    reg [7:0] out6409;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6409 = in0;
    end

    reg [7:0] out6410;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6410 = in0;
    end

    reg [7:0] out6411;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6411 = in0;
    end

    reg [7:0] out6412;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6412 = in0;
    end

    reg [7:0] out6413;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6413 = in0;
    end

    reg [7:0] out6414;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6414 = in0;
    end

    reg [7:0] out6415;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6415 = in0;
    end

    reg [7:0] out6416;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6416 = in0;
    end

    reg [7:0] out6417;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6417 = in0;
    end

    reg [7:0] out6418;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6418 = in0;
    end

    reg [7:0] out6419;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6419 = in0;
    end

    reg [7:0] out6420;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6420 = in0;
    end

    reg [7:0] out6421;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6421 = in0;
    end

    reg [7:0] out6422;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6422 = in0;
    end

    reg [7:0] out6423;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6423 = in0;
    end

    reg [7:0] out6424;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6424 = in0;
    end

    reg [7:0] out6425;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6425 = in0;
    end

    reg [7:0] out6426;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6426 = in0;
    end

    reg [7:0] out6427;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6427 = in0;
    end

    reg [7:0] out6428;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6428 = in0;
    end

    reg [7:0] out6429;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6429 = in0;
    end

    reg [7:0] out6430;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6430 = in0;
    end

    reg [7:0] out6431;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6431 = in0;
    end

    reg [7:0] out6432;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6432 = in0;
    end

    reg [7:0] out6433;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6433 = in0;
    end

    reg [7:0] out6434;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6434 = in0;
    end

    reg [7:0] out6435;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6435 = in0;
    end

    reg [7:0] out6436;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6436 = in0;
    end

    reg [7:0] out6437;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6437 = in0;
    end

    reg [7:0] out6438;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6438 = in0;
    end

    reg [7:0] out6439;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6439 = in0;
    end

    reg [7:0] out6440;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6440 = in0;
    end

    reg [7:0] out6441;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6441 = in0;
    end

    reg [7:0] out6442;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6442 = in0;
    end

    reg [7:0] out6443;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6443 = in0;
    end

    reg [7:0] out6444;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6444 = in0;
    end

    reg [7:0] out6445;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6445 = in0;
    end

    reg [7:0] out6446;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6446 = in0;
    end

    reg [7:0] out6447;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6447 = in0;
    end

    reg [7:0] out6448;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6448 = in0;
    end

    reg [7:0] out6449;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6449 = in0;
    end

    reg [7:0] out6450;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6450 = in0;
    end

    reg [7:0] out6451;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6451 = in0;
    end

    reg [7:0] out6452;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6452 = in0;
    end

    reg [7:0] out6453;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6453 = in0;
    end

    reg [7:0] out6454;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6454 = in0;
    end

    reg [7:0] out6455;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6455 = in0;
    end

    reg [7:0] out6456;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6456 = in0;
    end

    reg [7:0] out6457;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6457 = in0;
    end

    reg [7:0] out6458;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6458 = in0;
    end

    reg [7:0] out6459;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6459 = in0;
    end

    reg [7:0] out6460;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6460 = in0;
    end

    reg [7:0] out6461;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6461 = in0;
    end

    reg [7:0] out6462;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6462 = in0;
    end

    reg [7:0] out6463;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6463 = in0;
    end

    reg [7:0] out6464;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6464 = in0;
    end

    reg [7:0] out6465;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6465 = in0;
    end

    reg [7:0] out6466;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6466 = in0;
    end

    reg [7:0] out6467;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6467 = in0;
    end

    reg [7:0] out6468;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6468 = in0;
    end

    reg [7:0] out6469;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6469 = in0;
    end

    reg [7:0] out6470;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6470 = in0;
    end

    reg [7:0] out6471;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6471 = in0;
    end

    reg [7:0] out6472;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6472 = in0;
    end

    reg [7:0] out6473;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6473 = in0;
    end

    reg [7:0] out6474;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6474 = in0;
    end

    reg [7:0] out6475;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6475 = in0;
    end

    reg [7:0] out6476;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6476 = in0;
    end

    reg [7:0] out6477;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6477 = in0;
    end

    reg [7:0] out6478;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6478 = in0;
    end

    reg [7:0] out6479;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6479 = in0;
    end

    reg [7:0] out6480;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6480 = in0;
    end

    reg [7:0] out6481;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6481 = in0;
    end

    reg [7:0] out6482;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6482 = in0;
    end

    reg [7:0] out6483;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6483 = in0;
    end

    reg [7:0] out6484;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6484 = in0;
    end

    reg [7:0] out6485;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6485 = in0;
    end

    reg [7:0] out6486;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6486 = in0;
    end

    reg [7:0] out6487;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6487 = in0;
    end

    reg [7:0] out6488;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6488 = in0;
    end

    reg [7:0] out6489;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6489 = in0;
    end

    reg [7:0] out6490;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6490 = in0;
    end

    reg [7:0] out6491;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6491 = in0;
    end

    reg [7:0] out6492;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6492 = in0;
    end

    reg [7:0] out6493;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6493 = in0;
    end

    reg [7:0] out6494;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6494 = in0;
    end

    reg [7:0] out6495;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6495 = in0;
    end

    reg [7:0] out6496;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6496 = in0;
    end

    reg [7:0] out6497;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6497 = in0;
    end

    reg [7:0] out6498;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6498 = in0;
    end

    reg [7:0] out6499;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6499 = in0;
    end

    reg [7:0] out6500;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6500 = in0;
    end

    reg [7:0] out6501;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6501 = in0;
    end

    reg [7:0] out6502;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6502 = in0;
    end

    reg [7:0] out6503;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6503 = in0;
    end

    reg [7:0] out6504;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6504 = in0;
    end

    reg [7:0] out6505;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6505 = in0;
    end

    reg [7:0] out6506;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6506 = in0;
    end

    reg [7:0] out6507;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6507 = in0;
    end

    reg [7:0] out6508;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6508 = in0;
    end

    reg [7:0] out6509;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6509 = in0;
    end

    reg [7:0] out6510;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6510 = in0;
    end

    reg [7:0] out6511;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6511 = in0;
    end

    reg [7:0] out6512;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6512 = in0;
    end

    reg [7:0] out6513;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6513 = in0;
    end

    reg [7:0] out6514;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6514 = in0;
    end

    reg [7:0] out6515;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6515 = in0;
    end

    reg [7:0] out6516;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6516 = in0;
    end

    reg [7:0] out6517;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6517 = in0;
    end

    reg [7:0] out6518;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6518 = in0;
    end

    reg [7:0] out6519;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6519 = in0;
    end

    reg [7:0] out6520;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6520 = in0;
    end

    reg [7:0] out6521;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6521 = in0;
    end

    reg [7:0] out6522;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6522 = in0;
    end

    reg [7:0] out6523;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6523 = in0;
    end

    reg [7:0] out6524;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6524 = in0;
    end

    reg [7:0] out6525;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6525 = in0;
    end

    reg [7:0] out6526;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6526 = in0;
    end

    reg [7:0] out6527;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6527 = in0;
    end

    reg [7:0] out6528;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6528 = in0;
    end

    reg [7:0] out6529;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6529 = in0;
    end

    reg [7:0] out6530;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6530 = in0;
    end

    reg [7:0] out6531;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6531 = in0;
    end

    reg [7:0] out6532;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6532 = in0;
    end

    reg [7:0] out6533;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6533 = in0;
    end

    reg [7:0] out6534;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6534 = in0;
    end

    reg [7:0] out6535;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6535 = in0;
    end

    reg [7:0] out6536;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6536 = in0;
    end

    reg [7:0] out6537;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6537 = in0;
    end

    reg [7:0] out6538;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6538 = in0;
    end

    reg [7:0] out6539;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6539 = in0;
    end

    reg [7:0] out6540;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6540 = in0;
    end

    reg [7:0] out6541;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6541 = in0;
    end

    reg [7:0] out6542;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6542 = in0;
    end

    reg [7:0] out6543;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6543 = in0;
    end

    reg [7:0] out6544;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6544 = in0;
    end

    reg [7:0] out6545;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6545 = in0;
    end

    reg [7:0] out6546;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6546 = in0;
    end

    reg [7:0] out6547;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6547 = in0;
    end

    reg [7:0] out6548;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6548 = in0;
    end

    reg [7:0] out6549;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6549 = in0;
    end

    reg [7:0] out6550;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6550 = in0;
    end

    reg [7:0] out6551;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6551 = in0;
    end

    reg [7:0] out6552;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6552 = in0;
    end

    reg [7:0] out6553;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6553 = in0;
    end

    reg [7:0] out6554;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6554 = in0;
    end

    reg [7:0] out6555;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6555 = in0;
    end

    reg [7:0] out6556;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6556 = in0;
    end

    reg [7:0] out6557;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6557 = in0;
    end

    reg [7:0] out6558;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6558 = in0;
    end

    reg [7:0] out6559;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6559 = in0;
    end

    reg [7:0] out6560;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6560 = in0;
    end

    reg [7:0] out6561;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6561 = in0;
    end

    reg [7:0] out6562;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6562 = in0;
    end

    reg [7:0] out6563;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6563 = in0;
    end

    reg [7:0] out6564;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6564 = in0;
    end

    reg [7:0] out6565;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6565 = in0;
    end

    reg [7:0] out6566;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6566 = in0;
    end

    reg [7:0] out6567;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6567 = in0;
    end

    reg [7:0] out6568;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6568 = in0;
    end

    reg [7:0] out6569;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6569 = in0;
    end

    reg [7:0] out6570;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6570 = in0;
    end

    reg [7:0] out6571;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6571 = in0;
    end

    reg [7:0] out6572;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6572 = in0;
    end

    reg [7:0] out6573;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6573 = in0;
    end

    reg [7:0] out6574;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6574 = in0;
    end

    reg [7:0] out6575;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6575 = in0;
    end

    reg [7:0] out6576;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6576 = in0;
    end

    reg [7:0] out6577;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6577 = in0;
    end

    reg [7:0] out6578;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6578 = in0;
    end

    reg [7:0] out6579;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6579 = in0;
    end

    reg [7:0] out6580;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6580 = in0;
    end

    reg [7:0] out6581;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6581 = in0;
    end

    reg [7:0] out6582;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6582 = in0;
    end

    reg [7:0] out6583;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6583 = in0;
    end

    reg [7:0] out6584;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6584 = in0;
    end

    reg [7:0] out6585;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6585 = in0;
    end

    reg [7:0] out6586;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6586 = in0;
    end

    reg [7:0] out6587;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6587 = in0;
    end

    reg [7:0] out6588;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6588 = in0;
    end

    reg [7:0] out6589;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6589 = in0;
    end

    reg [7:0] out6590;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6590 = in0;
    end

    reg [7:0] out6591;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6591 = in0;
    end

    reg [7:0] out6592;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6592 = in0;
    end

    reg [7:0] out6593;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6593 = in0;
    end

    reg [7:0] out6594;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6594 = in0;
    end

    reg [7:0] out6595;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6595 = in0;
    end

    reg [7:0] out6596;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6596 = in0;
    end

    reg [7:0] out6597;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6597 = in0;
    end

    reg [7:0] out6598;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6598 = in0;
    end

    reg [7:0] out6599;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6599 = in0;
    end

    reg [7:0] out6600;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6600 = in0;
    end

    reg [7:0] out6601;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6601 = in0;
    end

    reg [7:0] out6602;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6602 = in0;
    end

    reg [7:0] out6603;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6603 = in0;
    end

    reg [7:0] out6604;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6604 = in0;
    end

    reg [7:0] out6605;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6605 = in0;
    end

    reg [7:0] out6606;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6606 = in0;
    end

    reg [7:0] out6607;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6607 = in0;
    end

    reg [7:0] out6608;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6608 = in0;
    end

    reg [7:0] out6609;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6609 = in0;
    end

    reg [7:0] out6610;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6610 = in0;
    end

    reg [7:0] out6611;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6611 = in0;
    end

    reg [7:0] out6612;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6612 = in0;
    end

    reg [7:0] out6613;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6613 = in0;
    end

    reg [7:0] out6614;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6614 = in0;
    end

    reg [7:0] out6615;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6615 = in0;
    end

    reg [7:0] out6616;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6616 = in0;
    end

    reg [7:0] out6617;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6617 = in0;
    end

    reg [7:0] out6618;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6618 = in0;
    end

    reg [7:0] out6619;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6619 = in0;
    end

    reg [7:0] out6620;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6620 = in0;
    end

    reg [7:0] out6621;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6621 = in0;
    end

    reg [7:0] out6622;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6622 = in0;
    end

    reg [7:0] out6623;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6623 = in0;
    end

    reg [7:0] out6624;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6624 = in0;
    end

    reg [7:0] out6625;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6625 = in0;
    end

    reg [7:0] out6626;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6626 = in0;
    end

    reg [7:0] out6627;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6627 = in0;
    end

    reg [7:0] out6628;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6628 = in0;
    end

    reg [7:0] out6629;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6629 = in0;
    end

    reg [7:0] out6630;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6630 = in0;
    end

    reg [7:0] out6631;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6631 = in0;
    end

    reg [7:0] out6632;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6632 = in0;
    end

    reg [7:0] out6633;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6633 = in0;
    end

    reg [7:0] out6634;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6634 = in0;
    end

    reg [7:0] out6635;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6635 = in0;
    end

    reg [7:0] out6636;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6636 = in0;
    end

    reg [7:0] out6637;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6637 = in0;
    end

    reg [7:0] out6638;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6638 = in0;
    end

    reg [7:0] out6639;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6639 = in0;
    end

    reg [7:0] out6640;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6640 = in0;
    end

    reg [7:0] out6641;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6641 = in0;
    end

    reg [7:0] out6642;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6642 = in0;
    end

    reg [7:0] out6643;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6643 = in0;
    end

    reg [7:0] out6644;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6644 = in0;
    end

    reg [7:0] out6645;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6645 = in0;
    end

    reg [7:0] out6646;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6646 = in0;
    end

    reg [7:0] out6647;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6647 = in0;
    end

    reg [7:0] out6648;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6648 = in0;
    end

    reg [7:0] out6649;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6649 = in0;
    end

    reg [7:0] out6650;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6650 = in0;
    end

    reg [7:0] out6651;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6651 = in0;
    end

    reg [7:0] out6652;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6652 = in0;
    end

    reg [7:0] out6653;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6653 = in0;
    end

    reg [7:0] out6654;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6654 = in0;
    end

    reg [7:0] out6655;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6655 = in0;
    end

    reg [7:0] out6656;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6656 = in0;
    end

    reg [7:0] out6657;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6657 = in0;
    end

    reg [7:0] out6658;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6658 = in0;
    end

    reg [7:0] out6659;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6659 = in0;
    end

    reg [7:0] out6660;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6660 = in0;
    end

    reg [7:0] out6661;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6661 = in0;
    end

    reg [7:0] out6662;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6662 = in0;
    end

    reg [7:0] out6663;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6663 = in0;
    end

    reg [7:0] out6664;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6664 = in0;
    end

    reg [7:0] out6665;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6665 = in0;
    end

    reg [7:0] out6666;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6666 = in0;
    end

    reg [7:0] out6667;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6667 = in0;
    end

    reg [7:0] out6668;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6668 = in0;
    end

    reg [7:0] out6669;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6669 = in0;
    end

    reg [7:0] out6670;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6670 = in0;
    end

    reg [7:0] out6671;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6671 = in0;
    end

    reg [7:0] out6672;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6672 = in0;
    end

    reg [7:0] out6673;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6673 = in0;
    end

    reg [7:0] out6674;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6674 = in0;
    end

    reg [7:0] out6675;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6675 = in0;
    end

    reg [7:0] out6676;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6676 = in0;
    end

    reg [7:0] out6677;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6677 = in0;
    end

    reg [7:0] out6678;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6678 = in0;
    end

    reg [7:0] out6679;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6679 = in0;
    end

    reg [7:0] out6680;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6680 = in0;
    end

    reg [7:0] out6681;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6681 = in0;
    end

    reg [7:0] out6682;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6682 = in0;
    end

    reg [7:0] out6683;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6683 = in0;
    end

    reg [7:0] out6684;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6684 = in0;
    end

    reg [7:0] out6685;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6685 = in0;
    end

    reg [7:0] out6686;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6686 = in0;
    end

    reg [7:0] out6687;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6687 = in0;
    end

    reg [7:0] out6688;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6688 = in0;
    end

    reg [7:0] out6689;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6689 = in0;
    end

    reg [7:0] out6690;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6690 = in0;
    end

    reg [7:0] out6691;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6691 = in0;
    end

    reg [7:0] out6692;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6692 = in0;
    end

    reg [7:0] out6693;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6693 = in0;
    end

    reg [7:0] out6694;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6694 = in0;
    end

    reg [7:0] out6695;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6695 = in0;
    end

    reg [7:0] out6696;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6696 = in0;
    end

    reg [7:0] out6697;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6697 = in0;
    end

    reg [7:0] out6698;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6698 = in0;
    end

    reg [7:0] out6699;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6699 = in0;
    end

    reg [7:0] out6700;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6700 = in0;
    end

    reg [7:0] out6701;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6701 = in0;
    end

    reg [7:0] out6702;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6702 = in0;
    end

    reg [7:0] out6703;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6703 = in0;
    end

    reg [7:0] out6704;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6704 = in0;
    end

    reg [7:0] out6705;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6705 = in0;
    end

    reg [7:0] out6706;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6706 = in0;
    end

    reg [7:0] out6707;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6707 = in0;
    end

    reg [7:0] out6708;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6708 = in0;
    end

    reg [7:0] out6709;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6709 = in0;
    end

    reg [7:0] out6710;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6710 = in0;
    end

    reg [7:0] out6711;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6711 = in0;
    end

    reg [7:0] out6712;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6712 = in0;
    end

    reg [7:0] out6713;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6713 = in0;
    end

    reg [7:0] out6714;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6714 = in0;
    end

    reg [7:0] out6715;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6715 = in0;
    end

    reg [7:0] out6716;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6716 = in0;
    end

    reg [7:0] out6717;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6717 = in0;
    end

    reg [7:0] out6718;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6718 = in0;
    end

    reg [7:0] out6719;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6719 = in0;
    end

    reg [7:0] out6720;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6720 = in0;
    end

    reg [7:0] out6721;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6721 = in0;
    end

    reg [7:0] out6722;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6722 = in0;
    end

    reg [7:0] out6723;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6723 = in0;
    end

    reg [7:0] out6724;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6724 = in0;
    end

    reg [7:0] out6725;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6725 = in0;
    end

    reg [7:0] out6726;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6726 = in0;
    end

    reg [7:0] out6727;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6727 = in0;
    end

    reg [7:0] out6728;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6728 = in0;
    end

    reg [7:0] out6729;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6729 = in0;
    end

    reg [7:0] out6730;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6730 = in0;
    end

    reg [7:0] out6731;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6731 = in0;
    end

    reg [7:0] out6732;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6732 = in0;
    end

    reg [7:0] out6733;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6733 = in0;
    end

    reg [7:0] out6734;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6734 = in0;
    end

    reg [7:0] out6735;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6735 = in0;
    end

    reg [7:0] out6736;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6736 = in0;
    end

    reg [7:0] out6737;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6737 = in0;
    end

    reg [7:0] out6738;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6738 = in0;
    end

    reg [7:0] out6739;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6739 = in0;
    end

    reg [7:0] out6740;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6740 = in0;
    end

    reg [7:0] out6741;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6741 = in0;
    end

    reg [7:0] out6742;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6742 = in0;
    end

    reg [7:0] out6743;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6743 = in0;
    end

    reg [7:0] out6744;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6744 = in0;
    end

    reg [7:0] out6745;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6745 = in0;
    end

    reg [7:0] out6746;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6746 = in0;
    end

    reg [7:0] out6747;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6747 = in0;
    end

    reg [7:0] out6748;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6748 = in0;
    end

    reg [7:0] out6749;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6749 = in0;
    end

    reg [7:0] out6750;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6750 = in0;
    end

    reg [7:0] out6751;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6751 = in0;
    end

    reg [7:0] out6752;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6752 = in0;
    end

    reg [7:0] out6753;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6753 = in0;
    end

    reg [7:0] out6754;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6754 = in0;
    end

    reg [7:0] out6755;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6755 = in0;
    end

    reg [7:0] out6756;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6756 = in0;
    end

    reg [7:0] out6757;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6757 = in0;
    end

    reg [7:0] out6758;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6758 = in0;
    end

    reg [7:0] out6759;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6759 = in0;
    end

    reg [7:0] out6760;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6760 = in0;
    end

    reg [7:0] out6761;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6761 = in0;
    end

    reg [7:0] out6762;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6762 = in0;
    end

    reg [7:0] out6763;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6763 = in0;
    end

    reg [7:0] out6764;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6764 = in0;
    end

    reg [7:0] out6765;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6765 = in0;
    end

    reg [7:0] out6766;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6766 = in0;
    end

    reg [7:0] out6767;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6767 = in0;
    end

    reg [7:0] out6768;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6768 = in0;
    end

    reg [7:0] out6769;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6769 = in0;
    end

    reg [7:0] out6770;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6770 = in0;
    end

    reg [7:0] out6771;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6771 = in0;
    end

    reg [7:0] out6772;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6772 = in0;
    end

    reg [7:0] out6773;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6773 = in0;
    end

    reg [7:0] out6774;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6774 = in0;
    end

    reg [7:0] out6775;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6775 = in0;
    end

    reg [7:0] out6776;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6776 = in0;
    end

    reg [7:0] out6777;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6777 = in0;
    end

    reg [7:0] out6778;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6778 = in0;
    end

    reg [7:0] out6779;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6779 = in0;
    end

    reg [7:0] out6780;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6780 = in0;
    end

    reg [7:0] out6781;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6781 = in0;
    end

    reg [7:0] out6782;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6782 = in0;
    end

    reg [7:0] out6783;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6783 = in0;
    end

    reg [7:0] out6784;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6784 = in0;
    end

    reg [7:0] out6785;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6785 = in0;
    end

    reg [7:0] out6786;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6786 = in0;
    end

    reg [7:0] out6787;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6787 = in0;
    end

    reg [7:0] out6788;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6788 = in0;
    end

    reg [7:0] out6789;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6789 = in0;
    end

    reg [7:0] out6790;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6790 = in0;
    end

    reg [7:0] out6791;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6791 = in0;
    end

    reg [7:0] out6792;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6792 = in0;
    end

    reg [7:0] out6793;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6793 = in0;
    end

    reg [7:0] out6794;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6794 = in0;
    end

    reg [7:0] out6795;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6795 = in0;
    end

    reg [7:0] out6796;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6796 = in0;
    end

    reg [7:0] out6797;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6797 = in0;
    end

    reg [7:0] out6798;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6798 = in0;
    end

    reg [7:0] out6799;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6799 = in0;
    end

    reg [7:0] out6800;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6800 = in0;
    end

    reg [7:0] out6801;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6801 = in0;
    end

    reg [7:0] out6802;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6802 = in0;
    end

    reg [7:0] out6803;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6803 = in0;
    end

    reg [7:0] out6804;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6804 = in0;
    end

    reg [7:0] out6805;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6805 = in0;
    end

    reg [7:0] out6806;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6806 = in0;
    end

    reg [7:0] out6807;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6807 = in0;
    end

    reg [7:0] out6808;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6808 = in0;
    end

    reg [7:0] out6809;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6809 = in0;
    end

    reg [7:0] out6810;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6810 = in0;
    end

    reg [7:0] out6811;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6811 = in0;
    end

    reg [7:0] out6812;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6812 = in0;
    end

    reg [7:0] out6813;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6813 = in0;
    end

    reg [7:0] out6814;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6814 = in0;
    end

    reg [7:0] out6815;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6815 = in0;
    end

    reg [7:0] out6816;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6816 = in0;
    end

    reg [7:0] out6817;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6817 = in0;
    end

    reg [7:0] out6818;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6818 = in0;
    end

    reg [7:0] out6819;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6819 = in0;
    end

    reg [7:0] out6820;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6820 = in0;
    end

    reg [7:0] out6821;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6821 = in0;
    end

    reg [7:0] out6822;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6822 = in0;
    end

    reg [7:0] out6823;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6823 = in0;
    end

    reg [7:0] out6824;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6824 = in0;
    end

    reg [7:0] out6825;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6825 = in0;
    end

    reg [7:0] out6826;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6826 = in0;
    end

    reg [7:0] out6827;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6827 = in0;
    end

    reg [7:0] out6828;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6828 = in0;
    end

    reg [7:0] out6829;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6829 = in0;
    end

    reg [7:0] out6830;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6830 = in0;
    end

    reg [7:0] out6831;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6831 = in0;
    end

    reg [7:0] out6832;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6832 = in0;
    end

    reg [7:0] out6833;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6833 = in0;
    end

    reg [7:0] out6834;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6834 = in0;
    end

    reg [7:0] out6835;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6835 = in0;
    end

    reg [7:0] out6836;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6836 = in0;
    end

    reg [7:0] out6837;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6837 = in0;
    end

    reg [7:0] out6838;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6838 = in0;
    end

    reg [7:0] out6839;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6839 = in0;
    end

    reg [7:0] out6840;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6840 = in0;
    end

    reg [7:0] out6841;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6841 = in0;
    end

    reg [7:0] out6842;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6842 = in0;
    end

    reg [7:0] out6843;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6843 = in0;
    end

    reg [7:0] out6844;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6844 = in0;
    end

    reg [7:0] out6845;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6845 = in0;
    end

    reg [7:0] out6846;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6846 = in0;
    end

    reg [7:0] out6847;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6847 = in0;
    end

    reg [7:0] out6848;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6848 = in0;
    end

    reg [7:0] out6849;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6849 = in0;
    end

    reg [7:0] out6850;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6850 = in0;
    end

    reg [7:0] out6851;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6851 = in0;
    end

    reg [7:0] out6852;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6852 = in0;
    end

    reg [7:0] out6853;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6853 = in0;
    end

    reg [7:0] out6854;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6854 = in0;
    end

    reg [7:0] out6855;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6855 = in0;
    end

    reg [7:0] out6856;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6856 = in0;
    end

    reg [7:0] out6857;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6857 = in0;
    end

    reg [7:0] out6858;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6858 = in0;
    end

    reg [7:0] out6859;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6859 = in0;
    end

    reg [7:0] out6860;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6860 = in0;
    end

    reg [7:0] out6861;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6861 = in0;
    end

    reg [7:0] out6862;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6862 = in0;
    end

    reg [7:0] out6863;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6863 = in0;
    end

    reg [7:0] out6864;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6864 = in0;
    end

    reg [7:0] out6865;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6865 = in0;
    end

    reg [7:0] out6866;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6866 = in0;
    end

    reg [7:0] out6867;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6867 = in0;
    end

    reg [7:0] out6868;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6868 = in0;
    end

    reg [7:0] out6869;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6869 = in0;
    end

    reg [7:0] out6870;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6870 = in0;
    end

    reg [7:0] out6871;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6871 = in0;
    end

    reg [7:0] out6872;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6872 = in0;
    end

    reg [7:0] out6873;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6873 = in0;
    end

    reg [7:0] out6874;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6874 = in0;
    end

    reg [7:0] out6875;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6875 = in0;
    end

    reg [7:0] out6876;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6876 = in0;
    end

    reg [7:0] out6877;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6877 = in0;
    end

    reg [7:0] out6878;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6878 = in0;
    end

    reg [7:0] out6879;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6879 = in0;
    end

    reg [7:0] out6880;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6880 = in0;
    end

    reg [7:0] out6881;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6881 = in0;
    end

    reg [7:0] out6882;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6882 = in0;
    end

    reg [7:0] out6883;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6883 = in0;
    end

    reg [7:0] out6884;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6884 = in0;
    end

    reg [7:0] out6885;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6885 = in0;
    end

    reg [7:0] out6886;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6886 = in0;
    end

    reg [7:0] out6887;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6887 = in0;
    end

    reg [7:0] out6888;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6888 = in0;
    end

    reg [7:0] out6889;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6889 = in0;
    end

    reg [7:0] out6890;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6890 = in0;
    end

    reg [7:0] out6891;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6891 = in0;
    end

    reg [7:0] out6892;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6892 = in0;
    end

    reg [7:0] out6893;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6893 = in0;
    end

    reg [7:0] out6894;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6894 = in0;
    end

    reg [7:0] out6895;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6895 = in0;
    end

    reg [7:0] out6896;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6896 = in0;
    end

    reg [7:0] out6897;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6897 = in0;
    end

    reg [7:0] out6898;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6898 = in0;
    end

    reg [7:0] out6899;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6899 = in0;
    end

    reg [7:0] out6900;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6900 = in0;
    end

    reg [7:0] out6901;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6901 = in0;
    end

    reg [7:0] out6902;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6902 = in0;
    end

    reg [7:0] out6903;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6903 = in0;
    end

    reg [7:0] out6904;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6904 = in0;
    end

    reg [7:0] out6905;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6905 = in0;
    end

    reg [7:0] out6906;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6906 = in0;
    end

    reg [7:0] out6907;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6907 = in0;
    end

    reg [7:0] out6908;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6908 = in0;
    end

    reg [7:0] out6909;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6909 = in0;
    end

    reg [7:0] out6910;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6910 = in0;
    end

    reg [7:0] out6911;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6911 = in0;
    end

    reg [7:0] out6912;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6912 = in0;
    end

    reg [7:0] out6913;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6913 = in0;
    end

    reg [7:0] out6914;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6914 = in0;
    end

    reg [7:0] out6915;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6915 = in0;
    end

    reg [7:0] out6916;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6916 = in0;
    end

    reg [7:0] out6917;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6917 = in0;
    end

    reg [7:0] out6918;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6918 = in0;
    end

    reg [7:0] out6919;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6919 = in0;
    end

    reg [7:0] out6920;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6920 = in0;
    end

    reg [7:0] out6921;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6921 = in0;
    end

    reg [7:0] out6922;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6922 = in0;
    end

    reg [7:0] out6923;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6923 = in0;
    end

    reg [7:0] out6924;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6924 = in0;
    end

    reg [7:0] out6925;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6925 = in0;
    end

    reg [7:0] out6926;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6926 = in0;
    end

    reg [7:0] out6927;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6927 = in0;
    end

    reg [7:0] out6928;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6928 = in0;
    end

    reg [7:0] out6929;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6929 = in0;
    end

    reg [7:0] out6930;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6930 = in0;
    end

    reg [7:0] out6931;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6931 = in0;
    end

    reg [7:0] out6932;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6932 = in0;
    end

    reg [7:0] out6933;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6933 = in0;
    end

    reg [7:0] out6934;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6934 = in0;
    end

    reg [7:0] out6935;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6935 = in0;
    end

    reg [7:0] out6936;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6936 = in0;
    end

    reg [7:0] out6937;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6937 = in0;
    end

    reg [7:0] out6938;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6938 = in0;
    end

    reg [7:0] out6939;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6939 = in0;
    end

    reg [7:0] out6940;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6940 = in0;
    end

    reg [7:0] out6941;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6941 = in0;
    end

    reg [7:0] out6942;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6942 = in0;
    end

    reg [7:0] out6943;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6943 = in0;
    end

    reg [7:0] out6944;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6944 = in0;
    end

    reg [7:0] out6945;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6945 = in0;
    end

    reg [7:0] out6946;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6946 = in0;
    end

    reg [7:0] out6947;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6947 = in0;
    end

    reg [7:0] out6948;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6948 = in0;
    end

    reg [7:0] out6949;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6949 = in0;
    end

    reg [7:0] out6950;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6950 = in0;
    end

    reg [7:0] out6951;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6951 = in0;
    end

    reg [7:0] out6952;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6952 = in0;
    end

    reg [7:0] out6953;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6953 = in0;
    end

    reg [7:0] out6954;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6954 = in0;
    end

    reg [7:0] out6955;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6955 = in0;
    end

    reg [7:0] out6956;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6956 = in0;
    end

    reg [7:0] out6957;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6957 = in0;
    end

    reg [7:0] out6958;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6958 = in0;
    end

    reg [7:0] out6959;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6959 = in0;
    end

    reg [7:0] out6960;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6960 = in0;
    end

    reg [7:0] out6961;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6961 = in0;
    end

    reg [7:0] out6962;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6962 = in0;
    end

    reg [7:0] out6963;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6963 = in0;
    end

    reg [7:0] out6964;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6964 = in0;
    end

    reg [7:0] out6965;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6965 = in0;
    end

    reg [7:0] out6966;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6966 = in0;
    end

    reg [7:0] out6967;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6967 = in0;
    end

    reg [7:0] out6968;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6968 = in0;
    end

    reg [7:0] out6969;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6969 = in0;
    end

    reg [7:0] out6970;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6970 = in0;
    end

    reg [7:0] out6971;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6971 = in0;
    end

    reg [7:0] out6972;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6972 = in0;
    end

    reg [7:0] out6973;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6973 = in0;
    end

    reg [7:0] out6974;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6974 = in0;
    end

    reg [7:0] out6975;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6975 = in0;
    end

    reg [7:0] out6976;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6976 = in0;
    end

    reg [7:0] out6977;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6977 = in0;
    end

    reg [7:0] out6978;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6978 = in0;
    end

    reg [7:0] out6979;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6979 = in0;
    end

    reg [7:0] out6980;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6980 = in0;
    end

    reg [7:0] out6981;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6981 = in0;
    end

    reg [7:0] out6982;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6982 = in0;
    end

    reg [7:0] out6983;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6983 = in0;
    end

    reg [7:0] out6984;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6984 = in0;
    end

    reg [7:0] out6985;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6985 = in0;
    end

    reg [7:0] out6986;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6986 = in0;
    end

    reg [7:0] out6987;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6987 = in0;
    end

    reg [7:0] out6988;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6988 = in0;
    end

    reg [7:0] out6989;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6989 = in0;
    end

    reg [7:0] out6990;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6990 = in0;
    end

    reg [7:0] out6991;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6991 = in0;
    end

    reg [7:0] out6992;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6992 = in0;
    end

    reg [7:0] out6993;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6993 = in0;
    end

    reg [7:0] out6994;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6994 = in0;
    end

    reg [7:0] out6995;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6995 = in0;
    end

    reg [7:0] out6996;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6996 = in0;
    end

    reg [7:0] out6997;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6997 = in0;
    end

    reg [7:0] out6998;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6998 = in0;
    end

    reg [7:0] out6999;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out6999 = in0;
    end

    reg [7:0] out7000;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7000 = in0;
    end

    reg [7:0] out7001;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7001 = in0;
    end

    reg [7:0] out7002;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7002 = in0;
    end

    reg [7:0] out7003;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7003 = in0;
    end

    reg [7:0] out7004;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7004 = in0;
    end

    reg [7:0] out7005;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7005 = in0;
    end

    reg [7:0] out7006;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7006 = in0;
    end

    reg [7:0] out7007;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7007 = in0;
    end

    reg [7:0] out7008;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7008 = in0;
    end

    reg [7:0] out7009;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7009 = in0;
    end

    reg [7:0] out7010;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7010 = in0;
    end

    reg [7:0] out7011;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7011 = in0;
    end

    reg [7:0] out7012;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7012 = in0;
    end

    reg [7:0] out7013;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7013 = in0;
    end

    reg [7:0] out7014;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7014 = in0;
    end

    reg [7:0] out7015;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7015 = in0;
    end

    reg [7:0] out7016;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7016 = in0;
    end

    reg [7:0] out7017;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7017 = in0;
    end

    reg [7:0] out7018;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7018 = in0;
    end

    reg [7:0] out7019;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7019 = in0;
    end

    reg [7:0] out7020;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7020 = in0;
    end

    reg [7:0] out7021;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7021 = in0;
    end

    reg [7:0] out7022;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7022 = in0;
    end

    reg [7:0] out7023;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7023 = in0;
    end

    reg [7:0] out7024;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7024 = in0;
    end

    reg [7:0] out7025;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7025 = in0;
    end

    reg [7:0] out7026;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7026 = in0;
    end

    reg [7:0] out7027;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7027 = in0;
    end

    reg [7:0] out7028;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7028 = in0;
    end

    reg [7:0] out7029;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7029 = in0;
    end

    reg [7:0] out7030;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7030 = in0;
    end

    reg [7:0] out7031;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7031 = in0;
    end

    reg [7:0] out7032;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7032 = in0;
    end

    reg [7:0] out7033;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7033 = in0;
    end

    reg [7:0] out7034;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7034 = in0;
    end

    reg [7:0] out7035;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7035 = in0;
    end

    reg [7:0] out7036;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7036 = in0;
    end

    reg [7:0] out7037;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7037 = in0;
    end

    reg [7:0] out7038;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7038 = in0;
    end

    reg [7:0] out7039;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7039 = in0;
    end

    reg [7:0] out7040;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7040 = in0;
    end

    reg [7:0] out7041;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7041 = in0;
    end

    reg [7:0] out7042;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7042 = in0;
    end

    reg [7:0] out7043;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7043 = in0;
    end

    reg [7:0] out7044;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7044 = in0;
    end

    reg [7:0] out7045;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7045 = in0;
    end

    reg [7:0] out7046;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7046 = in0;
    end

    reg [7:0] out7047;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7047 = in0;
    end

    reg [7:0] out7048;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7048 = in0;
    end

    reg [7:0] out7049;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7049 = in0;
    end

    reg [7:0] out7050;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7050 = in0;
    end

    reg [7:0] out7051;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7051 = in0;
    end

    reg [7:0] out7052;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7052 = in0;
    end

    reg [7:0] out7053;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7053 = in0;
    end

    reg [7:0] out7054;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7054 = in0;
    end

    reg [7:0] out7055;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7055 = in0;
    end

    reg [7:0] out7056;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7056 = in0;
    end

    reg [7:0] out7057;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7057 = in0;
    end

    reg [7:0] out7058;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7058 = in0;
    end

    reg [7:0] out7059;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7059 = in0;
    end

    reg [7:0] out7060;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7060 = in0;
    end

    reg [7:0] out7061;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7061 = in0;
    end

    reg [7:0] out7062;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7062 = in0;
    end

    reg [7:0] out7063;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7063 = in0;
    end

    reg [7:0] out7064;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7064 = in0;
    end

    reg [7:0] out7065;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7065 = in0;
    end

    reg [7:0] out7066;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7066 = in0;
    end

    reg [7:0] out7067;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7067 = in0;
    end

    reg [7:0] out7068;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7068 = in0;
    end

    reg [7:0] out7069;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7069 = in0;
    end

    reg [7:0] out7070;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7070 = in0;
    end

    reg [7:0] out7071;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7071 = in0;
    end

    reg [7:0] out7072;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7072 = in0;
    end

    reg [7:0] out7073;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7073 = in0;
    end

    reg [7:0] out7074;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7074 = in0;
    end

    reg [7:0] out7075;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7075 = in0;
    end

    reg [7:0] out7076;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7076 = in0;
    end

    reg [7:0] out7077;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7077 = in0;
    end

    reg [7:0] out7078;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7078 = in0;
    end

    reg [7:0] out7079;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7079 = in0;
    end

    reg [7:0] out7080;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7080 = in0;
    end

    reg [7:0] out7081;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7081 = in0;
    end

    reg [7:0] out7082;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7082 = in0;
    end

    reg [7:0] out7083;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7083 = in0;
    end

    reg [7:0] out7084;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7084 = in0;
    end

    reg [7:0] out7085;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7085 = in0;
    end

    reg [7:0] out7086;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7086 = in0;
    end

    reg [7:0] out7087;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7087 = in0;
    end

    reg [7:0] out7088;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7088 = in0;
    end

    reg [7:0] out7089;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7089 = in0;
    end

    reg [7:0] out7090;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7090 = in0;
    end

    reg [7:0] out7091;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7091 = in0;
    end

    reg [7:0] out7092;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7092 = in0;
    end

    reg [7:0] out7093;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7093 = in0;
    end

    reg [7:0] out7094;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7094 = in0;
    end

    reg [7:0] out7095;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7095 = in0;
    end

    reg [7:0] out7096;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7096 = in0;
    end

    reg [7:0] out7097;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7097 = in0;
    end

    reg [7:0] out7098;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7098 = in0;
    end

    reg [7:0] out7099;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7099 = in0;
    end

    reg [7:0] out7100;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7100 = in0;
    end

    reg [7:0] out7101;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7101 = in0;
    end

    reg [7:0] out7102;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7102 = in0;
    end

    reg [7:0] out7103;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7103 = in0;
    end

    reg [7:0] out7104;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7104 = in0;
    end

    reg [7:0] out7105;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7105 = in0;
    end

    reg [7:0] out7106;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7106 = in0;
    end

    reg [7:0] out7107;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7107 = in0;
    end

    reg [7:0] out7108;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7108 = in0;
    end

    reg [7:0] out7109;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7109 = in0;
    end

    reg [7:0] out7110;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7110 = in0;
    end

    reg [7:0] out7111;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7111 = in0;
    end

    reg [7:0] out7112;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7112 = in0;
    end

    reg [7:0] out7113;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7113 = in0;
    end

    reg [7:0] out7114;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7114 = in0;
    end

    reg [7:0] out7115;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7115 = in0;
    end

    reg [7:0] out7116;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7116 = in0;
    end

    reg [7:0] out7117;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7117 = in0;
    end

    reg [7:0] out7118;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7118 = in0;
    end

    reg [7:0] out7119;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7119 = in0;
    end

    reg [7:0] out7120;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7120 = in0;
    end

    reg [7:0] out7121;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7121 = in0;
    end

    reg [7:0] out7122;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7122 = in0;
    end

    reg [7:0] out7123;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7123 = in0;
    end

    reg [7:0] out7124;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7124 = in0;
    end

    reg [7:0] out7125;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7125 = in0;
    end

    reg [7:0] out7126;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7126 = in0;
    end

    reg [7:0] out7127;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7127 = in0;
    end

    reg [7:0] out7128;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7128 = in0;
    end

    reg [7:0] out7129;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7129 = in0;
    end

    reg [7:0] out7130;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7130 = in0;
    end

    reg [7:0] out7131;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7131 = in0;
    end

    reg [7:0] out7132;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7132 = in0;
    end

    reg [7:0] out7133;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7133 = in0;
    end

    reg [7:0] out7134;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7134 = in0;
    end

    reg [7:0] out7135;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7135 = in0;
    end

    reg [7:0] out7136;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7136 = in0;
    end

    reg [7:0] out7137;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7137 = in0;
    end

    reg [7:0] out7138;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7138 = in0;
    end

    reg [7:0] out7139;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7139 = in0;
    end

    reg [7:0] out7140;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7140 = in0;
    end

    reg [7:0] out7141;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7141 = in0;
    end

    reg [7:0] out7142;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7142 = in0;
    end

    reg [7:0] out7143;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7143 = in0;
    end

    reg [7:0] out7144;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7144 = in0;
    end

    reg [7:0] out7145;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7145 = in0;
    end

    reg [7:0] out7146;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7146 = in0;
    end

    reg [7:0] out7147;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7147 = in0;
    end

    reg [7:0] out7148;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7148 = in0;
    end

    reg [7:0] out7149;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7149 = in0;
    end

    reg [7:0] out7150;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7150 = in0;
    end

    reg [7:0] out7151;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7151 = in0;
    end

    reg [7:0] out7152;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7152 = in0;
    end

    reg [7:0] out7153;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7153 = in0;
    end

    reg [7:0] out7154;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7154 = in0;
    end

    reg [7:0] out7155;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7155 = in0;
    end

    reg [7:0] out7156;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7156 = in0;
    end

    reg [7:0] out7157;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7157 = in0;
    end

    reg [7:0] out7158;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7158 = in0;
    end

    reg [7:0] out7159;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7159 = in0;
    end

    reg [7:0] out7160;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7160 = in0;
    end

    reg [7:0] out7161;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7161 = in0;
    end

    reg [7:0] out7162;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7162 = in0;
    end

    reg [7:0] out7163;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7163 = in0;
    end

    reg [7:0] out7164;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7164 = in0;
    end

    reg [7:0] out7165;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7165 = in0;
    end

    reg [7:0] out7166;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7166 = in0;
    end

    reg [7:0] out7167;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7167 = in0;
    end

    reg [7:0] out7168;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7168 = in0;
    end

    reg [7:0] out7169;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7169 = in0;
    end

    reg [7:0] out7170;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7170 = in0;
    end

    reg [7:0] out7171;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7171 = in0;
    end

    reg [7:0] out7172;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7172 = in0;
    end

    reg [7:0] out7173;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7173 = in0;
    end

    reg [7:0] out7174;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7174 = in0;
    end

    reg [7:0] out7175;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7175 = in0;
    end

    reg [7:0] out7176;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7176 = in0;
    end

    reg [7:0] out7177;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7177 = in0;
    end

    reg [7:0] out7178;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7178 = in0;
    end

    reg [7:0] out7179;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7179 = in0;
    end

    reg [7:0] out7180;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7180 = in0;
    end

    reg [7:0] out7181;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7181 = in0;
    end

    reg [7:0] out7182;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7182 = in0;
    end

    reg [7:0] out7183;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7183 = in0;
    end

    reg [7:0] out7184;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7184 = in0;
    end

    reg [7:0] out7185;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7185 = in0;
    end

    reg [7:0] out7186;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7186 = in0;
    end

    reg [7:0] out7187;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7187 = in0;
    end

    reg [7:0] out7188;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7188 = in0;
    end

    reg [7:0] out7189;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7189 = in0;
    end

    reg [7:0] out7190;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7190 = in0;
    end

    reg [7:0] out7191;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7191 = in0;
    end

    reg [7:0] out7192;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7192 = in0;
    end

    reg [7:0] out7193;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7193 = in0;
    end

    reg [7:0] out7194;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7194 = in0;
    end

    reg [7:0] out7195;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7195 = in0;
    end

    reg [7:0] out7196;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7196 = in0;
    end

    reg [7:0] out7197;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7197 = in0;
    end

    reg [7:0] out7198;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7198 = in0;
    end

    reg [7:0] out7199;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7199 = in0;
    end

    reg [7:0] out7200;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7200 = in0;
    end

    reg [7:0] out7201;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7201 = in0;
    end

    reg [7:0] out7202;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7202 = in0;
    end

    reg [7:0] out7203;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7203 = in0;
    end

    reg [7:0] out7204;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7204 = in0;
    end

    reg [7:0] out7205;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7205 = in0;
    end

    reg [7:0] out7206;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7206 = in0;
    end

    reg [7:0] out7207;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7207 = in0;
    end

    reg [7:0] out7208;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7208 = in0;
    end

    reg [7:0] out7209;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7209 = in0;
    end

    reg [7:0] out7210;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7210 = in0;
    end

    reg [7:0] out7211;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7211 = in0;
    end

    reg [7:0] out7212;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7212 = in0;
    end

    reg [7:0] out7213;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7213 = in0;
    end

    reg [7:0] out7214;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7214 = in0;
    end

    reg [7:0] out7215;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7215 = in0;
    end

    reg [7:0] out7216;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7216 = in0;
    end

    reg [7:0] out7217;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7217 = in0;
    end

    reg [7:0] out7218;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7218 = in0;
    end

    reg [7:0] out7219;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7219 = in0;
    end

    reg [7:0] out7220;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7220 = in0;
    end

    reg [7:0] out7221;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7221 = in0;
    end

    reg [7:0] out7222;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7222 = in0;
    end

    reg [7:0] out7223;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7223 = in0;
    end

    reg [7:0] out7224;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7224 = in0;
    end

    reg [7:0] out7225;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7225 = in0;
    end

    reg [7:0] out7226;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7226 = in0;
    end

    reg [7:0] out7227;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7227 = in0;
    end

    reg [7:0] out7228;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7228 = in0;
    end

    reg [7:0] out7229;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7229 = in0;
    end

    reg [7:0] out7230;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7230 = in0;
    end

    reg [7:0] out7231;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7231 = in0;
    end

    reg [7:0] out7232;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7232 = in0;
    end

    reg [7:0] out7233;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7233 = in0;
    end

    reg [7:0] out7234;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7234 = in0;
    end

    reg [7:0] out7235;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7235 = in0;
    end

    reg [7:0] out7236;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7236 = in0;
    end

    reg [7:0] out7237;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7237 = in0;
    end

    reg [7:0] out7238;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7238 = in0;
    end

    reg [7:0] out7239;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7239 = in0;
    end

    reg [7:0] out7240;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7240 = in0;
    end

    reg [7:0] out7241;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7241 = in0;
    end

    reg [7:0] out7242;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7242 = in0;
    end

    reg [7:0] out7243;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7243 = in0;
    end

    reg [7:0] out7244;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7244 = in0;
    end

    reg [7:0] out7245;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7245 = in0;
    end

    reg [7:0] out7246;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7246 = in0;
    end

    reg [7:0] out7247;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7247 = in0;
    end

    reg [7:0] out7248;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7248 = in0;
    end

    reg [7:0] out7249;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7249 = in0;
    end

    reg [7:0] out7250;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7250 = in0;
    end

    reg [7:0] out7251;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7251 = in0;
    end

    reg [7:0] out7252;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7252 = in0;
    end

    reg [7:0] out7253;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7253 = in0;
    end

    reg [7:0] out7254;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7254 = in0;
    end

    reg [7:0] out7255;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7255 = in0;
    end

    reg [7:0] out7256;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7256 = in0;
    end

    reg [7:0] out7257;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7257 = in0;
    end

    reg [7:0] out7258;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7258 = in0;
    end

    reg [7:0] out7259;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7259 = in0;
    end

    reg [7:0] out7260;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7260 = in0;
    end

    reg [7:0] out7261;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7261 = in0;
    end

    reg [7:0] out7262;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7262 = in0;
    end

    reg [7:0] out7263;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7263 = in0;
    end

    reg [7:0] out7264;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7264 = in0;
    end

    reg [7:0] out7265;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7265 = in0;
    end

    reg [7:0] out7266;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7266 = in0;
    end

    reg [7:0] out7267;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7267 = in0;
    end

    reg [7:0] out7268;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7268 = in0;
    end

    reg [7:0] out7269;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7269 = in0;
    end

    reg [7:0] out7270;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7270 = in0;
    end

    reg [7:0] out7271;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7271 = in0;
    end

    reg [7:0] out7272;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7272 = in0;
    end

    reg [7:0] out7273;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7273 = in0;
    end

    reg [7:0] out7274;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7274 = in0;
    end

    reg [7:0] out7275;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7275 = in0;
    end

    reg [7:0] out7276;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7276 = in0;
    end

    reg [7:0] out7277;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7277 = in0;
    end

    reg [7:0] out7278;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7278 = in0;
    end

    reg [7:0] out7279;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7279 = in0;
    end

    reg [7:0] out7280;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7280 = in0;
    end

    reg [7:0] out7281;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7281 = in0;
    end

    reg [7:0] out7282;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7282 = in0;
    end

    reg [7:0] out7283;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7283 = in0;
    end

    reg [7:0] out7284;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7284 = in0;
    end

    reg [7:0] out7285;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7285 = in0;
    end

    reg [7:0] out7286;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7286 = in0;
    end

    reg [7:0] out7287;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7287 = in0;
    end

    reg [7:0] out7288;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7288 = in0;
    end

    reg [7:0] out7289;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7289 = in0;
    end

    reg [7:0] out7290;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7290 = in0;
    end

    reg [7:0] out7291;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7291 = in0;
    end

    reg [7:0] out7292;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7292 = in0;
    end

    reg [7:0] out7293;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7293 = in0;
    end

    reg [7:0] out7294;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7294 = in0;
    end

    reg [7:0] out7295;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7295 = in0;
    end

    reg [7:0] out7296;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7296 = in0;
    end

    reg [7:0] out7297;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7297 = in0;
    end

    reg [7:0] out7298;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7298 = in0;
    end

    reg [7:0] out7299;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7299 = in0;
    end

    reg [7:0] out7300;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7300 = in0;
    end

    reg [7:0] out7301;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7301 = in0;
    end

    reg [7:0] out7302;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7302 = in0;
    end

    reg [7:0] out7303;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7303 = in0;
    end

    reg [7:0] out7304;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7304 = in0;
    end

    reg [7:0] out7305;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7305 = in0;
    end

    reg [7:0] out7306;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7306 = in0;
    end

    reg [7:0] out7307;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7307 = in0;
    end

    reg [7:0] out7308;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7308 = in0;
    end

    reg [7:0] out7309;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7309 = in0;
    end

    reg [7:0] out7310;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7310 = in0;
    end

    reg [7:0] out7311;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7311 = in0;
    end

    reg [7:0] out7312;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7312 = in0;
    end

    reg [7:0] out7313;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7313 = in0;
    end

    reg [7:0] out7314;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7314 = in0;
    end

    reg [7:0] out7315;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7315 = in0;
    end

    reg [7:0] out7316;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7316 = in0;
    end

    reg [7:0] out7317;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7317 = in0;
    end

    reg [7:0] out7318;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7318 = in0;
    end

    reg [7:0] out7319;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7319 = in0;
    end

    reg [7:0] out7320;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7320 = in0;
    end

    reg [7:0] out7321;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7321 = in0;
    end

    reg [7:0] out7322;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7322 = in0;
    end

    reg [7:0] out7323;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7323 = in0;
    end

    reg [7:0] out7324;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7324 = in0;
    end

    reg [7:0] out7325;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7325 = in0;
    end

    reg [7:0] out7326;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7326 = in0;
    end

    reg [7:0] out7327;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7327 = in0;
    end

    reg [7:0] out7328;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7328 = in0;
    end

    reg [7:0] out7329;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7329 = in0;
    end

    reg [7:0] out7330;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7330 = in0;
    end

    reg [7:0] out7331;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7331 = in0;
    end

    reg [7:0] out7332;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7332 = in0;
    end

    reg [7:0] out7333;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7333 = in0;
    end

    reg [7:0] out7334;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7334 = in0;
    end

    reg [7:0] out7335;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7335 = in0;
    end

    reg [7:0] out7336;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7336 = in0;
    end

    reg [7:0] out7337;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7337 = in0;
    end

    reg [7:0] out7338;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7338 = in0;
    end

    reg [7:0] out7339;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7339 = in0;
    end

    reg [7:0] out7340;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7340 = in0;
    end

    reg [7:0] out7341;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7341 = in0;
    end

    reg [7:0] out7342;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7342 = in0;
    end

    reg [7:0] out7343;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7343 = in0;
    end

    reg [7:0] out7344;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7344 = in0;
    end

    reg [7:0] out7345;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7345 = in0;
    end

    reg [7:0] out7346;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7346 = in0;
    end

    reg [7:0] out7347;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7347 = in0;
    end

    reg [7:0] out7348;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7348 = in0;
    end

    reg [7:0] out7349;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7349 = in0;
    end

    reg [7:0] out7350;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7350 = in0;
    end

    reg [7:0] out7351;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7351 = in0;
    end

    reg [7:0] out7352;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7352 = in0;
    end

    reg [7:0] out7353;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7353 = in0;
    end

    reg [7:0] out7354;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7354 = in0;
    end

    reg [7:0] out7355;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7355 = in0;
    end

    reg [7:0] out7356;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7356 = in0;
    end

    reg [7:0] out7357;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7357 = in0;
    end

    reg [7:0] out7358;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7358 = in0;
    end

    reg [7:0] out7359;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7359 = in0;
    end

    reg [7:0] out7360;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7360 = in0;
    end

    reg [7:0] out7361;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7361 = in0;
    end

    reg [7:0] out7362;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7362 = in0;
    end

    reg [7:0] out7363;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7363 = in0;
    end

    reg [7:0] out7364;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7364 = in0;
    end

    reg [7:0] out7365;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7365 = in0;
    end

    reg [7:0] out7366;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7366 = in0;
    end

    reg [7:0] out7367;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7367 = in0;
    end

    reg [7:0] out7368;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7368 = in0;
    end

    reg [7:0] out7369;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7369 = in0;
    end

    reg [7:0] out7370;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7370 = in0;
    end

    reg [7:0] out7371;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7371 = in0;
    end

    reg [7:0] out7372;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7372 = in0;
    end

    reg [7:0] out7373;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7373 = in0;
    end

    reg [7:0] out7374;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7374 = in0;
    end

    reg [7:0] out7375;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7375 = in0;
    end

    reg [7:0] out7376;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7376 = in0;
    end

    reg [7:0] out7377;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7377 = in0;
    end

    reg [7:0] out7378;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7378 = in0;
    end

    reg [7:0] out7379;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7379 = in0;
    end

    reg [7:0] out7380;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7380 = in0;
    end

    reg [7:0] out7381;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7381 = in0;
    end

    reg [7:0] out7382;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7382 = in0;
    end

    reg [7:0] out7383;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7383 = in0;
    end

    reg [7:0] out7384;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7384 = in0;
    end

    reg [7:0] out7385;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7385 = in0;
    end

    reg [7:0] out7386;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7386 = in0;
    end

    reg [7:0] out7387;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7387 = in0;
    end

    reg [7:0] out7388;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7388 = in0;
    end

    reg [7:0] out7389;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7389 = in0;
    end

    reg [7:0] out7390;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7390 = in0;
    end

    reg [7:0] out7391;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7391 = in0;
    end

    reg [7:0] out7392;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7392 = in0;
    end

    reg [7:0] out7393;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7393 = in0;
    end

    reg [7:0] out7394;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7394 = in0;
    end

    reg [7:0] out7395;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7395 = in0;
    end

    reg [7:0] out7396;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7396 = in0;
    end

    reg [7:0] out7397;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7397 = in0;
    end

    reg [7:0] out7398;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7398 = in0;
    end

    reg [7:0] out7399;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7399 = in0;
    end

    reg [7:0] out7400;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7400 = in0;
    end

    reg [7:0] out7401;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7401 = in0;
    end

    reg [7:0] out7402;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7402 = in0;
    end

    reg [7:0] out7403;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7403 = in0;
    end

    reg [7:0] out7404;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7404 = in0;
    end

    reg [7:0] out7405;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7405 = in0;
    end

    reg [7:0] out7406;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7406 = in0;
    end

    reg [7:0] out7407;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7407 = in0;
    end

    reg [7:0] out7408;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7408 = in0;
    end

    reg [7:0] out7409;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7409 = in0;
    end

    reg [7:0] out7410;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7410 = in0;
    end

    reg [7:0] out7411;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7411 = in0;
    end

    reg [7:0] out7412;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7412 = in0;
    end

    reg [7:0] out7413;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7413 = in0;
    end

    reg [7:0] out7414;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7414 = in0;
    end

    reg [7:0] out7415;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7415 = in0;
    end

    reg [7:0] out7416;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7416 = in0;
    end

    reg [7:0] out7417;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7417 = in0;
    end

    reg [7:0] out7418;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7418 = in0;
    end

    reg [7:0] out7419;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7419 = in0;
    end

    reg [7:0] out7420;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7420 = in0;
    end

    reg [7:0] out7421;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7421 = in0;
    end

    reg [7:0] out7422;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7422 = in0;
    end

    reg [7:0] out7423;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7423 = in0;
    end

    reg [7:0] out7424;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7424 = in0;
    end

    reg [7:0] out7425;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7425 = in0;
    end

    reg [7:0] out7426;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7426 = in0;
    end

    reg [7:0] out7427;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7427 = in0;
    end

    reg [7:0] out7428;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7428 = in0;
    end

    reg [7:0] out7429;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7429 = in0;
    end

    reg [7:0] out7430;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7430 = in0;
    end

    reg [7:0] out7431;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7431 = in0;
    end

    reg [7:0] out7432;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7432 = in0;
    end

    reg [7:0] out7433;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7433 = in0;
    end

    reg [7:0] out7434;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7434 = in0;
    end

    reg [7:0] out7435;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7435 = in0;
    end

    reg [7:0] out7436;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7436 = in0;
    end

    reg [7:0] out7437;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7437 = in0;
    end

    reg [7:0] out7438;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7438 = in0;
    end

    reg [7:0] out7439;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7439 = in0;
    end

    reg [7:0] out7440;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7440 = in0;
    end

    reg [7:0] out7441;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7441 = in0;
    end

    reg [7:0] out7442;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7442 = in0;
    end

    reg [7:0] out7443;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7443 = in0;
    end

    reg [7:0] out7444;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7444 = in0;
    end

    reg [7:0] out7445;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7445 = in0;
    end

    reg [7:0] out7446;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7446 = in0;
    end

    reg [7:0] out7447;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7447 = in0;
    end

    reg [7:0] out7448;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7448 = in0;
    end

    reg [7:0] out7449;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7449 = in0;
    end

    reg [7:0] out7450;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7450 = in0;
    end

    reg [7:0] out7451;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7451 = in0;
    end

    reg [7:0] out7452;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7452 = in0;
    end

    reg [7:0] out7453;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7453 = in0;
    end

    reg [7:0] out7454;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7454 = in0;
    end

    reg [7:0] out7455;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7455 = in0;
    end

    reg [7:0] out7456;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7456 = in0;
    end

    reg [7:0] out7457;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7457 = in0;
    end

    reg [7:0] out7458;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7458 = in0;
    end

    reg [7:0] out7459;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7459 = in0;
    end

    reg [7:0] out7460;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7460 = in0;
    end

    reg [7:0] out7461;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7461 = in0;
    end

    reg [7:0] out7462;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7462 = in0;
    end

    reg [7:0] out7463;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7463 = in0;
    end

    reg [7:0] out7464;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7464 = in0;
    end

    reg [7:0] out7465;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7465 = in0;
    end

    reg [7:0] out7466;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7466 = in0;
    end

    reg [7:0] out7467;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7467 = in0;
    end

    reg [7:0] out7468;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7468 = in0;
    end

    reg [7:0] out7469;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7469 = in0;
    end

    reg [7:0] out7470;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7470 = in0;
    end

    reg [7:0] out7471;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7471 = in0;
    end

    reg [7:0] out7472;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7472 = in0;
    end

    reg [7:0] out7473;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7473 = in0;
    end

    reg [7:0] out7474;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7474 = in0;
    end

    reg [7:0] out7475;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7475 = in0;
    end

    reg [7:0] out7476;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7476 = in0;
    end

    reg [7:0] out7477;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7477 = in0;
    end

    reg [7:0] out7478;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7478 = in0;
    end

    reg [7:0] out7479;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7479 = in0;
    end

    reg [7:0] out7480;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7480 = in0;
    end

    reg [7:0] out7481;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7481 = in0;
    end

    reg [7:0] out7482;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7482 = in0;
    end

    reg [7:0] out7483;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7483 = in0;
    end

    reg [7:0] out7484;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7484 = in0;
    end

    reg [7:0] out7485;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7485 = in0;
    end

    reg [7:0] out7486;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7486 = in0;
    end

    reg [7:0] out7487;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7487 = in0;
    end

    reg [7:0] out7488;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7488 = in0;
    end

    reg [7:0] out7489;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7489 = in0;
    end

    reg [7:0] out7490;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7490 = in0;
    end

    reg [7:0] out7491;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7491 = in0;
    end

    reg [7:0] out7492;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7492 = in0;
    end

    reg [7:0] out7493;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7493 = in0;
    end

    reg [7:0] out7494;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7494 = in0;
    end

    reg [7:0] out7495;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7495 = in0;
    end

    reg [7:0] out7496;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7496 = in0;
    end

    reg [7:0] out7497;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7497 = in0;
    end

    reg [7:0] out7498;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7498 = in0;
    end

    reg [7:0] out7499;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7499 = in0;
    end

    reg [7:0] out7500;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7500 = in0;
    end

    reg [7:0] out7501;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7501 = in0;
    end

    reg [7:0] out7502;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7502 = in0;
    end

    reg [7:0] out7503;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7503 = in0;
    end

    reg [7:0] out7504;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7504 = in0;
    end

    reg [7:0] out7505;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7505 = in0;
    end

    reg [7:0] out7506;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7506 = in0;
    end

    reg [7:0] out7507;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7507 = in0;
    end

    reg [7:0] out7508;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7508 = in0;
    end

    reg [7:0] out7509;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7509 = in0;
    end

    reg [7:0] out7510;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7510 = in0;
    end

    reg [7:0] out7511;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7511 = in0;
    end

    reg [7:0] out7512;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7512 = in0;
    end

    reg [7:0] out7513;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7513 = in0;
    end

    reg [7:0] out7514;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7514 = in0;
    end

    reg [7:0] out7515;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7515 = in0;
    end

    reg [7:0] out7516;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7516 = in0;
    end

    reg [7:0] out7517;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7517 = in0;
    end

    reg [7:0] out7518;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7518 = in0;
    end

    reg [7:0] out7519;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7519 = in0;
    end

    reg [7:0] out7520;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7520 = in0;
    end

    reg [7:0] out7521;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7521 = in0;
    end

    reg [7:0] out7522;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7522 = in0;
    end

    reg [7:0] out7523;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7523 = in0;
    end

    reg [7:0] out7524;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7524 = in0;
    end

    reg [7:0] out7525;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7525 = in0;
    end

    reg [7:0] out7526;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7526 = in0;
    end

    reg [7:0] out7527;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7527 = in0;
    end

    reg [7:0] out7528;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7528 = in0;
    end

    reg [7:0] out7529;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7529 = in0;
    end

    reg [7:0] out7530;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7530 = in0;
    end

    reg [7:0] out7531;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7531 = in0;
    end

    reg [7:0] out7532;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7532 = in0;
    end

    reg [7:0] out7533;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7533 = in0;
    end

    reg [7:0] out7534;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7534 = in0;
    end

    reg [7:0] out7535;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7535 = in0;
    end

    reg [7:0] out7536;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7536 = in0;
    end

    reg [7:0] out7537;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7537 = in0;
    end

    reg [7:0] out7538;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7538 = in0;
    end

    reg [7:0] out7539;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7539 = in0;
    end

    reg [7:0] out7540;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7540 = in0;
    end

    reg [7:0] out7541;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7541 = in0;
    end

    reg [7:0] out7542;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7542 = in0;
    end

    reg [7:0] out7543;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7543 = in0;
    end

    reg [7:0] out7544;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7544 = in0;
    end

    reg [7:0] out7545;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7545 = in0;
    end

    reg [7:0] out7546;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7546 = in0;
    end

    reg [7:0] out7547;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7547 = in0;
    end

    reg [7:0] out7548;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7548 = in0;
    end

    reg [7:0] out7549;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7549 = in0;
    end

    reg [7:0] out7550;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7550 = in0;
    end

    reg [7:0] out7551;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7551 = in0;
    end

    reg [7:0] out7552;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7552 = in0;
    end

    reg [7:0] out7553;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7553 = in0;
    end

    reg [7:0] out7554;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7554 = in0;
    end

    reg [7:0] out7555;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7555 = in0;
    end

    reg [7:0] out7556;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7556 = in0;
    end

    reg [7:0] out7557;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7557 = in0;
    end

    reg [7:0] out7558;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7558 = in0;
    end

    reg [7:0] out7559;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7559 = in0;
    end

    reg [7:0] out7560;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7560 = in0;
    end

    reg [7:0] out7561;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7561 = in0;
    end

    reg [7:0] out7562;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7562 = in0;
    end

    reg [7:0] out7563;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7563 = in0;
    end

    reg [7:0] out7564;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7564 = in0;
    end

    reg [7:0] out7565;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7565 = in0;
    end

    reg [7:0] out7566;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7566 = in0;
    end

    reg [7:0] out7567;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7567 = in0;
    end

    reg [7:0] out7568;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7568 = in0;
    end

    reg [7:0] out7569;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7569 = in0;
    end

    reg [7:0] out7570;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7570 = in0;
    end

    reg [7:0] out7571;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7571 = in0;
    end

    reg [7:0] out7572;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7572 = in0;
    end

    reg [7:0] out7573;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7573 = in0;
    end

    reg [7:0] out7574;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7574 = in0;
    end

    reg [7:0] out7575;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7575 = in0;
    end

    reg [7:0] out7576;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7576 = in0;
    end

    reg [7:0] out7577;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7577 = in0;
    end

    reg [7:0] out7578;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7578 = in0;
    end

    reg [7:0] out7579;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7579 = in0;
    end

    reg [7:0] out7580;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7580 = in0;
    end

    reg [7:0] out7581;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7581 = in0;
    end

    reg [7:0] out7582;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7582 = in0;
    end

    reg [7:0] out7583;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7583 = in0;
    end

    reg [7:0] out7584;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7584 = in0;
    end

    reg [7:0] out7585;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7585 = in0;
    end

    reg [7:0] out7586;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7586 = in0;
    end

    reg [7:0] out7587;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7587 = in0;
    end

    reg [7:0] out7588;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7588 = in0;
    end

    reg [7:0] out7589;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7589 = in0;
    end

    reg [7:0] out7590;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7590 = in0;
    end

    reg [7:0] out7591;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7591 = in0;
    end

    reg [7:0] out7592;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7592 = in0;
    end

    reg [7:0] out7593;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7593 = in0;
    end

    reg [7:0] out7594;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7594 = in0;
    end

    reg [7:0] out7595;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7595 = in0;
    end

    reg [7:0] out7596;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7596 = in0;
    end

    reg [7:0] out7597;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7597 = in0;
    end

    reg [7:0] out7598;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7598 = in0;
    end

    reg [7:0] out7599;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7599 = in0;
    end

    reg [7:0] out7600;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7600 = in0;
    end

    reg [7:0] out7601;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7601 = in0;
    end

    reg [7:0] out7602;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7602 = in0;
    end

    reg [7:0] out7603;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7603 = in0;
    end

    reg [7:0] out7604;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7604 = in0;
    end

    reg [7:0] out7605;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7605 = in0;
    end

    reg [7:0] out7606;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7606 = in0;
    end

    reg [7:0] out7607;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7607 = in0;
    end

    reg [7:0] out7608;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7608 = in0;
    end

    reg [7:0] out7609;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7609 = in0;
    end

    reg [7:0] out7610;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7610 = in0;
    end

    reg [7:0] out7611;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7611 = in0;
    end

    reg [7:0] out7612;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7612 = in0;
    end

    reg [7:0] out7613;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7613 = in0;
    end

    reg [7:0] out7614;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7614 = in0;
    end

    reg [7:0] out7615;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7615 = in0;
    end

    reg [7:0] out7616;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7616 = in0;
    end

    reg [7:0] out7617;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7617 = in0;
    end

    reg [7:0] out7618;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7618 = in0;
    end

    reg [7:0] out7619;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7619 = in0;
    end

    reg [7:0] out7620;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7620 = in0;
    end

    reg [7:0] out7621;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7621 = in0;
    end

    reg [7:0] out7622;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7622 = in0;
    end

    reg [7:0] out7623;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7623 = in0;
    end

    reg [7:0] out7624;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7624 = in0;
    end

    reg [7:0] out7625;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7625 = in0;
    end

    reg [7:0] out7626;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7626 = in0;
    end

    reg [7:0] out7627;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7627 = in0;
    end

    reg [7:0] out7628;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7628 = in0;
    end

    reg [7:0] out7629;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7629 = in0;
    end

    reg [7:0] out7630;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7630 = in0;
    end

    reg [7:0] out7631;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7631 = in0;
    end

    reg [7:0] out7632;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7632 = in0;
    end

    reg [7:0] out7633;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7633 = in0;
    end

    reg [7:0] out7634;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7634 = in0;
    end

    reg [7:0] out7635;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7635 = in0;
    end

    reg [7:0] out7636;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7636 = in0;
    end

    reg [7:0] out7637;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7637 = in0;
    end

    reg [7:0] out7638;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7638 = in0;
    end

    reg [7:0] out7639;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7639 = in0;
    end

    reg [7:0] out7640;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7640 = in0;
    end

    reg [7:0] out7641;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7641 = in0;
    end

    reg [7:0] out7642;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7642 = in0;
    end

    reg [7:0] out7643;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7643 = in0;
    end

    reg [7:0] out7644;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7644 = in0;
    end

    reg [7:0] out7645;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7645 = in0;
    end

    reg [7:0] out7646;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7646 = in0;
    end

    reg [7:0] out7647;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7647 = in0;
    end

    reg [7:0] out7648;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7648 = in0;
    end

    reg [7:0] out7649;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7649 = in0;
    end

    reg [7:0] out7650;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7650 = in0;
    end

    reg [7:0] out7651;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7651 = in0;
    end

    reg [7:0] out7652;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7652 = in0;
    end

    reg [7:0] out7653;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7653 = in0;
    end

    reg [7:0] out7654;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7654 = in0;
    end

    reg [7:0] out7655;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7655 = in0;
    end

    reg [7:0] out7656;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7656 = in0;
    end

    reg [7:0] out7657;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7657 = in0;
    end

    reg [7:0] out7658;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7658 = in0;
    end

    reg [7:0] out7659;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7659 = in0;
    end

    reg [7:0] out7660;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7660 = in0;
    end

    reg [7:0] out7661;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7661 = in0;
    end

    reg [7:0] out7662;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7662 = in0;
    end

    reg [7:0] out7663;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7663 = in0;
    end

    reg [7:0] out7664;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7664 = in0;
    end

    reg [7:0] out7665;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7665 = in0;
    end

    reg [7:0] out7666;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7666 = in0;
    end

    reg [7:0] out7667;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7667 = in0;
    end

    reg [7:0] out7668;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7668 = in0;
    end

    reg [7:0] out7669;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7669 = in0;
    end

    reg [7:0] out7670;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7670 = in0;
    end

    reg [7:0] out7671;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7671 = in0;
    end

    reg [7:0] out7672;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7672 = in0;
    end

    reg [7:0] out7673;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7673 = in0;
    end

    reg [7:0] out7674;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7674 = in0;
    end

    reg [7:0] out7675;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7675 = in0;
    end

    reg [7:0] out7676;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7676 = in0;
    end

    reg [7:0] out7677;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7677 = in0;
    end

    reg [7:0] out7678;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7678 = in0;
    end

    reg [7:0] out7679;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7679 = in0;
    end

    reg [7:0] out7680;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7680 = in0;
    end

    reg [7:0] out7681;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7681 = in0;
    end

    reg [7:0] out7682;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7682 = in0;
    end

    reg [7:0] out7683;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7683 = in0;
    end

    reg [7:0] out7684;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7684 = in0;
    end

    reg [7:0] out7685;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7685 = in0;
    end

    reg [7:0] out7686;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7686 = in0;
    end

    reg [7:0] out7687;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7687 = in0;
    end

    reg [7:0] out7688;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7688 = in0;
    end

    reg [7:0] out7689;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7689 = in0;
    end

    reg [7:0] out7690;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7690 = in0;
    end

    reg [7:0] out7691;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7691 = in0;
    end

    reg [7:0] out7692;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7692 = in0;
    end

    reg [7:0] out7693;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7693 = in0;
    end

    reg [7:0] out7694;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7694 = in0;
    end

    reg [7:0] out7695;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7695 = in0;
    end

    reg [7:0] out7696;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7696 = in0;
    end

    reg [7:0] out7697;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7697 = in0;
    end

    reg [7:0] out7698;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7698 = in0;
    end

    reg [7:0] out7699;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7699 = in0;
    end

    reg [7:0] out7700;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7700 = in0;
    end

    reg [7:0] out7701;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7701 = in0;
    end

    reg [7:0] out7702;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7702 = in0;
    end

    reg [7:0] out7703;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7703 = in0;
    end

    reg [7:0] out7704;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7704 = in0;
    end

    reg [7:0] out7705;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7705 = in0;
    end

    reg [7:0] out7706;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7706 = in0;
    end

    reg [7:0] out7707;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7707 = in0;
    end

    reg [7:0] out7708;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7708 = in0;
    end

    reg [7:0] out7709;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7709 = in0;
    end

    reg [7:0] out7710;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7710 = in0;
    end

    reg [7:0] out7711;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7711 = in0;
    end

    reg [7:0] out7712;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7712 = in0;
    end

    reg [7:0] out7713;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7713 = in0;
    end

    reg [7:0] out7714;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7714 = in0;
    end

    reg [7:0] out7715;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7715 = in0;
    end

    reg [7:0] out7716;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7716 = in0;
    end

    reg [7:0] out7717;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7717 = in0;
    end

    reg [7:0] out7718;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7718 = in0;
    end

    reg [7:0] out7719;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7719 = in0;
    end

    reg [7:0] out7720;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7720 = in0;
    end

    reg [7:0] out7721;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7721 = in0;
    end

    reg [7:0] out7722;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7722 = in0;
    end

    reg [7:0] out7723;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7723 = in0;
    end

    reg [7:0] out7724;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7724 = in0;
    end

    reg [7:0] out7725;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7725 = in0;
    end

    reg [7:0] out7726;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7726 = in0;
    end

    reg [7:0] out7727;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7727 = in0;
    end

    reg [7:0] out7728;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7728 = in0;
    end

    reg [7:0] out7729;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7729 = in0;
    end

    reg [7:0] out7730;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7730 = in0;
    end

    reg [7:0] out7731;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7731 = in0;
    end

    reg [7:0] out7732;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7732 = in0;
    end

    reg [7:0] out7733;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7733 = in0;
    end

    reg [7:0] out7734;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7734 = in0;
    end

    reg [7:0] out7735;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7735 = in0;
    end

    reg [7:0] out7736;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7736 = in0;
    end

    reg [7:0] out7737;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7737 = in0;
    end

    reg [7:0] out7738;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7738 = in0;
    end

    reg [7:0] out7739;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7739 = in0;
    end

    reg [7:0] out7740;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7740 = in0;
    end

    reg [7:0] out7741;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7741 = in0;
    end

    reg [7:0] out7742;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7742 = in0;
    end

    reg [7:0] out7743;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7743 = in0;
    end

    reg [7:0] out7744;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7744 = in0;
    end

    reg [7:0] out7745;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7745 = in0;
    end

    reg [7:0] out7746;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7746 = in0;
    end

    reg [7:0] out7747;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7747 = in0;
    end

    reg [7:0] out7748;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7748 = in0;
    end

    reg [7:0] out7749;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7749 = in0;
    end

    reg [7:0] out7750;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7750 = in0;
    end

    reg [7:0] out7751;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7751 = in0;
    end

    reg [7:0] out7752;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7752 = in0;
    end

    reg [7:0] out7753;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7753 = in0;
    end

    reg [7:0] out7754;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7754 = in0;
    end

    reg [7:0] out7755;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7755 = in0;
    end

    reg [7:0] out7756;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7756 = in0;
    end

    reg [7:0] out7757;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7757 = in0;
    end

    reg [7:0] out7758;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7758 = in0;
    end

    reg [7:0] out7759;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7759 = in0;
    end

    reg [7:0] out7760;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7760 = in0;
    end

    reg [7:0] out7761;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7761 = in0;
    end

    reg [7:0] out7762;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7762 = in0;
    end

    reg [7:0] out7763;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7763 = in0;
    end

    reg [7:0] out7764;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7764 = in0;
    end

    reg [7:0] out7765;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7765 = in0;
    end

    reg [7:0] out7766;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7766 = in0;
    end

    reg [7:0] out7767;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7767 = in0;
    end

    reg [7:0] out7768;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7768 = in0;
    end

    reg [7:0] out7769;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7769 = in0;
    end

    reg [7:0] out7770;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7770 = in0;
    end

    reg [7:0] out7771;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7771 = in0;
    end

    reg [7:0] out7772;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7772 = in0;
    end

    reg [7:0] out7773;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7773 = in0;
    end

    reg [7:0] out7774;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7774 = in0;
    end

    reg [7:0] out7775;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7775 = in0;
    end

    reg [7:0] out7776;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7776 = in0;
    end

    reg [7:0] out7777;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7777 = in0;
    end

    reg [7:0] out7778;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7778 = in0;
    end

    reg [7:0] out7779;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7779 = in0;
    end

    reg [7:0] out7780;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7780 = in0;
    end

    reg [7:0] out7781;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7781 = in0;
    end

    reg [7:0] out7782;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7782 = in0;
    end

    reg [7:0] out7783;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7783 = in0;
    end

    reg [7:0] out7784;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7784 = in0;
    end

    reg [7:0] out7785;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7785 = in0;
    end

    reg [7:0] out7786;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7786 = in0;
    end

    reg [7:0] out7787;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7787 = in0;
    end

    reg [7:0] out7788;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7788 = in0;
    end

    reg [7:0] out7789;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7789 = in0;
    end

    reg [7:0] out7790;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7790 = in0;
    end

    reg [7:0] out7791;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7791 = in0;
    end

    reg [7:0] out7792;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7792 = in0;
    end

    reg [7:0] out7793;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7793 = in0;
    end

    reg [7:0] out7794;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7794 = in0;
    end

    reg [7:0] out7795;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7795 = in0;
    end

    reg [7:0] out7796;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7796 = in0;
    end

    reg [7:0] out7797;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7797 = in0;
    end

    reg [7:0] out7798;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7798 = in0;
    end

    reg [7:0] out7799;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7799 = in0;
    end

    reg [7:0] out7800;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7800 = in0;
    end

    reg [7:0] out7801;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7801 = in0;
    end

    reg [7:0] out7802;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7802 = in0;
    end

    reg [7:0] out7803;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7803 = in0;
    end

    reg [7:0] out7804;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7804 = in0;
    end

    reg [7:0] out7805;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7805 = in0;
    end

    reg [7:0] out7806;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7806 = in0;
    end

    reg [7:0] out7807;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7807 = in0;
    end

    reg [7:0] out7808;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7808 = in0;
    end

    reg [7:0] out7809;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7809 = in0;
    end

    reg [7:0] out7810;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7810 = in0;
    end

    reg [7:0] out7811;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7811 = in0;
    end

    reg [7:0] out7812;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7812 = in0;
    end

    reg [7:0] out7813;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7813 = in0;
    end

    reg [7:0] out7814;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7814 = in0;
    end

    reg [7:0] out7815;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7815 = in0;
    end

    reg [7:0] out7816;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7816 = in0;
    end

    reg [7:0] out7817;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7817 = in0;
    end

    reg [7:0] out7818;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7818 = in0;
    end

    reg [7:0] out7819;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7819 = in0;
    end

    reg [7:0] out7820;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7820 = in0;
    end

    reg [7:0] out7821;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7821 = in0;
    end

    reg [7:0] out7822;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7822 = in0;
    end

    reg [7:0] out7823;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7823 = in0;
    end

    reg [7:0] out7824;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7824 = in0;
    end

    reg [7:0] out7825;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7825 = in0;
    end

    reg [7:0] out7826;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7826 = in0;
    end

    reg [7:0] out7827;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7827 = in0;
    end

    reg [7:0] out7828;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7828 = in0;
    end

    reg [7:0] out7829;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7829 = in0;
    end

    reg [7:0] out7830;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7830 = in0;
    end

    reg [7:0] out7831;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7831 = in0;
    end

    reg [7:0] out7832;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7832 = in0;
    end

    reg [7:0] out7833;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7833 = in0;
    end

    reg [7:0] out7834;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7834 = in0;
    end

    reg [7:0] out7835;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7835 = in0;
    end

    reg [7:0] out7836;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7836 = in0;
    end

    reg [7:0] out7837;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7837 = in0;
    end

    reg [7:0] out7838;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7838 = in0;
    end

    reg [7:0] out7839;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7839 = in0;
    end

    reg [7:0] out7840;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7840 = in0;
    end

    reg [7:0] out7841;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7841 = in0;
    end

    reg [7:0] out7842;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7842 = in0;
    end

    reg [7:0] out7843;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7843 = in0;
    end

    reg [7:0] out7844;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7844 = in0;
    end

    reg [7:0] out7845;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7845 = in0;
    end

    reg [7:0] out7846;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7846 = in0;
    end

    reg [7:0] out7847;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7847 = in0;
    end

    reg [7:0] out7848;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7848 = in0;
    end

    reg [7:0] out7849;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7849 = in0;
    end

    reg [7:0] out7850;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7850 = in0;
    end

    reg [7:0] out7851;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7851 = in0;
    end

    reg [7:0] out7852;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7852 = in0;
    end

    reg [7:0] out7853;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7853 = in0;
    end

    reg [7:0] out7854;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7854 = in0;
    end

    reg [7:0] out7855;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7855 = in0;
    end

    reg [7:0] out7856;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7856 = in0;
    end

    reg [7:0] out7857;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7857 = in0;
    end

    reg [7:0] out7858;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7858 = in0;
    end

    reg [7:0] out7859;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7859 = in0;
    end

    reg [7:0] out7860;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7860 = in0;
    end

    reg [7:0] out7861;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7861 = in0;
    end

    reg [7:0] out7862;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7862 = in0;
    end

    reg [7:0] out7863;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7863 = in0;
    end

    reg [7:0] out7864;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7864 = in0;
    end

    reg [7:0] out7865;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7865 = in0;
    end

    reg [7:0] out7866;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7866 = in0;
    end

    reg [7:0] out7867;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7867 = in0;
    end

    reg [7:0] out7868;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7868 = in0;
    end

    reg [7:0] out7869;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7869 = in0;
    end

    reg [7:0] out7870;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7870 = in0;
    end

    reg [7:0] out7871;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7871 = in0;
    end

    reg [7:0] out7872;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7872 = in0;
    end

    reg [7:0] out7873;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7873 = in0;
    end

    reg [7:0] out7874;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7874 = in0;
    end

    reg [7:0] out7875;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7875 = in0;
    end

    reg [7:0] out7876;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7876 = in0;
    end

    reg [7:0] out7877;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7877 = in0;
    end

    reg [7:0] out7878;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7878 = in0;
    end

    reg [7:0] out7879;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7879 = in0;
    end

    reg [7:0] out7880;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7880 = in0;
    end

    reg [7:0] out7881;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7881 = in0;
    end

    reg [7:0] out7882;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7882 = in0;
    end

    reg [7:0] out7883;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7883 = in0;
    end

    reg [7:0] out7884;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7884 = in0;
    end

    reg [7:0] out7885;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7885 = in0;
    end

    reg [7:0] out7886;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7886 = in0;
    end

    reg [7:0] out7887;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7887 = in0;
    end

    reg [7:0] out7888;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7888 = in0;
    end

    reg [7:0] out7889;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7889 = in0;
    end

    reg [7:0] out7890;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7890 = in0;
    end

    reg [7:0] out7891;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7891 = in0;
    end

    reg [7:0] out7892;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7892 = in0;
    end

    reg [7:0] out7893;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7893 = in0;
    end

    reg [7:0] out7894;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7894 = in0;
    end

    reg [7:0] out7895;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7895 = in0;
    end

    reg [7:0] out7896;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7896 = in0;
    end

    reg [7:0] out7897;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7897 = in0;
    end

    reg [7:0] out7898;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7898 = in0;
    end

    reg [7:0] out7899;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7899 = in0;
    end

    reg [7:0] out7900;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7900 = in0;
    end

    reg [7:0] out7901;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7901 = in0;
    end

    reg [7:0] out7902;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7902 = in0;
    end

    reg [7:0] out7903;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7903 = in0;
    end

    reg [7:0] out7904;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7904 = in0;
    end

    reg [7:0] out7905;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7905 = in0;
    end

    reg [7:0] out7906;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7906 = in0;
    end

    reg [7:0] out7907;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7907 = in0;
    end

    reg [7:0] out7908;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7908 = in0;
    end

    reg [7:0] out7909;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7909 = in0;
    end

    reg [7:0] out7910;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7910 = in0;
    end

    reg [7:0] out7911;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7911 = in0;
    end

    reg [7:0] out7912;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7912 = in0;
    end

    reg [7:0] out7913;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7913 = in0;
    end

    reg [7:0] out7914;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7914 = in0;
    end

    reg [7:0] out7915;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7915 = in0;
    end

    reg [7:0] out7916;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7916 = in0;
    end

    reg [7:0] out7917;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7917 = in0;
    end

    reg [7:0] out7918;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7918 = in0;
    end

    reg [7:0] out7919;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7919 = in0;
    end

    reg [7:0] out7920;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7920 = in0;
    end

    reg [7:0] out7921;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7921 = in0;
    end

    reg [7:0] out7922;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7922 = in0;
    end

    reg [7:0] out7923;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7923 = in0;
    end

    reg [7:0] out7924;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7924 = in0;
    end

    reg [7:0] out7925;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7925 = in0;
    end

    reg [7:0] out7926;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7926 = in0;
    end

    reg [7:0] out7927;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7927 = in0;
    end

    reg [7:0] out7928;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7928 = in0;
    end

    reg [7:0] out7929;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7929 = in0;
    end

    reg [7:0] out7930;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7930 = in0;
    end

    reg [7:0] out7931;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7931 = in0;
    end

    reg [7:0] out7932;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7932 = in0;
    end

    reg [7:0] out7933;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7933 = in0;
    end

    reg [7:0] out7934;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7934 = in0;
    end

    reg [7:0] out7935;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7935 = in0;
    end

    reg [7:0] out7936;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7936 = in0;
    end

    reg [7:0] out7937;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7937 = in0;
    end

    reg [7:0] out7938;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7938 = in0;
    end

    reg [7:0] out7939;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7939 = in0;
    end

    reg [7:0] out7940;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7940 = in0;
    end

    reg [7:0] out7941;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7941 = in0;
    end

    reg [7:0] out7942;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7942 = in0;
    end

    reg [7:0] out7943;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7943 = in0;
    end

    reg [7:0] out7944;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7944 = in0;
    end

    reg [7:0] out7945;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7945 = in0;
    end

    reg [7:0] out7946;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7946 = in0;
    end

    reg [7:0] out7947;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7947 = in0;
    end

    reg [7:0] out7948;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7948 = in0;
    end

    reg [7:0] out7949;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7949 = in0;
    end

    reg [7:0] out7950;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7950 = in0;
    end

    reg [7:0] out7951;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7951 = in0;
    end

    reg [7:0] out7952;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7952 = in0;
    end

    reg [7:0] out7953;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7953 = in0;
    end

    reg [7:0] out7954;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7954 = in0;
    end

    reg [7:0] out7955;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7955 = in0;
    end

    reg [7:0] out7956;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7956 = in0;
    end

    reg [7:0] out7957;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7957 = in0;
    end

    reg [7:0] out7958;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7958 = in0;
    end

    reg [7:0] out7959;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7959 = in0;
    end

    reg [7:0] out7960;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7960 = in0;
    end

    reg [7:0] out7961;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7961 = in0;
    end

    reg [7:0] out7962;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7962 = in0;
    end

    reg [7:0] out7963;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7963 = in0;
    end

    reg [7:0] out7964;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7964 = in0;
    end

    reg [7:0] out7965;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7965 = in0;
    end

    reg [7:0] out7966;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7966 = in0;
    end

    reg [7:0] out7967;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7967 = in0;
    end

    reg [7:0] out7968;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7968 = in0;
    end

    reg [7:0] out7969;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7969 = in0;
    end

    reg [7:0] out7970;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7970 = in0;
    end

    reg [7:0] out7971;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7971 = in0;
    end

    reg [7:0] out7972;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7972 = in0;
    end

    reg [7:0] out7973;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7973 = in0;
    end

    reg [7:0] out7974;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7974 = in0;
    end

    reg [7:0] out7975;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7975 = in0;
    end

    reg [7:0] out7976;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7976 = in0;
    end

    reg [7:0] out7977;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7977 = in0;
    end

    reg [7:0] out7978;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7978 = in0;
    end

    reg [7:0] out7979;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7979 = in0;
    end

    reg [7:0] out7980;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7980 = in0;
    end

    reg [7:0] out7981;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7981 = in0;
    end

    reg [7:0] out7982;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7982 = in0;
    end

    reg [7:0] out7983;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7983 = in0;
    end

    reg [7:0] out7984;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7984 = in0;
    end

    reg [7:0] out7985;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7985 = in0;
    end

    reg [7:0] out7986;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7986 = in0;
    end

    reg [7:0] out7987;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7987 = in0;
    end

    reg [7:0] out7988;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7988 = in0;
    end

    reg [7:0] out7989;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7989 = in0;
    end

    reg [7:0] out7990;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7990 = in0;
    end

    reg [7:0] out7991;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7991 = in0;
    end

    reg [7:0] out7992;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7992 = in0;
    end

    reg [7:0] out7993;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7993 = in0;
    end

    reg [7:0] out7994;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7994 = in0;
    end

    reg [7:0] out7995;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7995 = in0;
    end

    reg [7:0] out7996;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7996 = in0;
    end

    reg [7:0] out7997;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7997 = in0;
    end

    reg [7:0] out7998;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7998 = in0;
    end

    reg [7:0] out7999;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out7999 = in0;
    end

    reg [7:0] out8000;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8000 = in0;
    end

    reg [7:0] out8001;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8001 = in0;
    end

    reg [7:0] out8002;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8002 = in0;
    end

    reg [7:0] out8003;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8003 = in0;
    end

    reg [7:0] out8004;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8004 = in0;
    end

    reg [7:0] out8005;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8005 = in0;
    end

    reg [7:0] out8006;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8006 = in0;
    end

    reg [7:0] out8007;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8007 = in0;
    end

    reg [7:0] out8008;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8008 = in0;
    end

    reg [7:0] out8009;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8009 = in0;
    end

    reg [7:0] out8010;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8010 = in0;
    end

    reg [7:0] out8011;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8011 = in0;
    end

    reg [7:0] out8012;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8012 = in0;
    end

    reg [7:0] out8013;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8013 = in0;
    end

    reg [7:0] out8014;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8014 = in0;
    end

    reg [7:0] out8015;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8015 = in0;
    end

    reg [7:0] out8016;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8016 = in0;
    end

    reg [7:0] out8017;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8017 = in0;
    end

    reg [7:0] out8018;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8018 = in0;
    end

    reg [7:0] out8019;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8019 = in0;
    end

    reg [7:0] out8020;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8020 = in0;
    end

    reg [7:0] out8021;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8021 = in0;
    end

    reg [7:0] out8022;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8022 = in0;
    end

    reg [7:0] out8023;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8023 = in0;
    end

    reg [7:0] out8024;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8024 = in0;
    end

    reg [7:0] out8025;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8025 = in0;
    end

    reg [7:0] out8026;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8026 = in0;
    end

    reg [7:0] out8027;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8027 = in0;
    end

    reg [7:0] out8028;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8028 = in0;
    end

    reg [7:0] out8029;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8029 = in0;
    end

    reg [7:0] out8030;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8030 = in0;
    end

    reg [7:0] out8031;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8031 = in0;
    end

    reg [7:0] out8032;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8032 = in0;
    end

    reg [7:0] out8033;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8033 = in0;
    end

    reg [7:0] out8034;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8034 = in0;
    end

    reg [7:0] out8035;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8035 = in0;
    end

    reg [7:0] out8036;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8036 = in0;
    end

    reg [7:0] out8037;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8037 = in0;
    end

    reg [7:0] out8038;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8038 = in0;
    end

    reg [7:0] out8039;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8039 = in0;
    end

    reg [7:0] out8040;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8040 = in0;
    end

    reg [7:0] out8041;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8041 = in0;
    end

    reg [7:0] out8042;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8042 = in0;
    end

    reg [7:0] out8043;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8043 = in0;
    end

    reg [7:0] out8044;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8044 = in0;
    end

    reg [7:0] out8045;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8045 = in0;
    end

    reg [7:0] out8046;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8046 = in0;
    end

    reg [7:0] out8047;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8047 = in0;
    end

    reg [7:0] out8048;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8048 = in0;
    end

    reg [7:0] out8049;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8049 = in0;
    end

    reg [7:0] out8050;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8050 = in0;
    end

    reg [7:0] out8051;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8051 = in0;
    end

    reg [7:0] out8052;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8052 = in0;
    end

    reg [7:0] out8053;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8053 = in0;
    end

    reg [7:0] out8054;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8054 = in0;
    end

    reg [7:0] out8055;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8055 = in0;
    end

    reg [7:0] out8056;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8056 = in0;
    end

    reg [7:0] out8057;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8057 = in0;
    end

    reg [7:0] out8058;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8058 = in0;
    end

    reg [7:0] out8059;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8059 = in0;
    end

    reg [7:0] out8060;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8060 = in0;
    end

    reg [7:0] out8061;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8061 = in0;
    end

    reg [7:0] out8062;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8062 = in0;
    end

    reg [7:0] out8063;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8063 = in0;
    end

    reg [7:0] out8064;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8064 = in0;
    end

    reg [7:0] out8065;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8065 = in0;
    end

    reg [7:0] out8066;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8066 = in0;
    end

    reg [7:0] out8067;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8067 = in0;
    end

    reg [7:0] out8068;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8068 = in0;
    end

    reg [7:0] out8069;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8069 = in0;
    end

    reg [7:0] out8070;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8070 = in0;
    end

    reg [7:0] out8071;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8071 = in0;
    end

    reg [7:0] out8072;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8072 = in0;
    end

    reg [7:0] out8073;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8073 = in0;
    end

    reg [7:0] out8074;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8074 = in0;
    end

    reg [7:0] out8075;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8075 = in0;
    end

    reg [7:0] out8076;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8076 = in0;
    end

    reg [7:0] out8077;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8077 = in0;
    end

    reg [7:0] out8078;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8078 = in0;
    end

    reg [7:0] out8079;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8079 = in0;
    end

    reg [7:0] out8080;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8080 = in0;
    end

    reg [7:0] out8081;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8081 = in0;
    end

    reg [7:0] out8082;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8082 = in0;
    end

    reg [7:0] out8083;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8083 = in0;
    end

    reg [7:0] out8084;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8084 = in0;
    end

    reg [7:0] out8085;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8085 = in0;
    end

    reg [7:0] out8086;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8086 = in0;
    end

    reg [7:0] out8087;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8087 = in0;
    end

    reg [7:0] out8088;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8088 = in0;
    end

    reg [7:0] out8089;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8089 = in0;
    end

    reg [7:0] out8090;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8090 = in0;
    end

    reg [7:0] out8091;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8091 = in0;
    end

    reg [7:0] out8092;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8092 = in0;
    end

    reg [7:0] out8093;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8093 = in0;
    end

    reg [7:0] out8094;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8094 = in0;
    end

    reg [7:0] out8095;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8095 = in0;
    end

    reg [7:0] out8096;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8096 = in0;
    end

    reg [7:0] out8097;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8097 = in0;
    end

    reg [7:0] out8098;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8098 = in0;
    end

    reg [7:0] out8099;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8099 = in0;
    end

    reg [7:0] out8100;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8100 = in0;
    end

    reg [7:0] out8101;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8101 = in0;
    end

    reg [7:0] out8102;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8102 = in0;
    end

    reg [7:0] out8103;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8103 = in0;
    end

    reg [7:0] out8104;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8104 = in0;
    end

    reg [7:0] out8105;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8105 = in0;
    end

    reg [7:0] out8106;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8106 = in0;
    end

    reg [7:0] out8107;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8107 = in0;
    end

    reg [7:0] out8108;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8108 = in0;
    end

    reg [7:0] out8109;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8109 = in0;
    end

    reg [7:0] out8110;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8110 = in0;
    end

    reg [7:0] out8111;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8111 = in0;
    end

    reg [7:0] out8112;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8112 = in0;
    end

    reg [7:0] out8113;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8113 = in0;
    end

    reg [7:0] out8114;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8114 = in0;
    end

    reg [7:0] out8115;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8115 = in0;
    end

    reg [7:0] out8116;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8116 = in0;
    end

    reg [7:0] out8117;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8117 = in0;
    end

    reg [7:0] out8118;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8118 = in0;
    end

    reg [7:0] out8119;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8119 = in0;
    end

    reg [7:0] out8120;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8120 = in0;
    end

    reg [7:0] out8121;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8121 = in0;
    end

    reg [7:0] out8122;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8122 = in0;
    end

    reg [7:0] out8123;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8123 = in0;
    end

    reg [7:0] out8124;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8124 = in0;
    end

    reg [7:0] out8125;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8125 = in0;
    end

    reg [7:0] out8126;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8126 = in0;
    end

    reg [7:0] out8127;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8127 = in0;
    end

    reg [7:0] out8128;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8128 = in0;
    end

    reg [7:0] out8129;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8129 = in0;
    end

    reg [7:0] out8130;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8130 = in0;
    end

    reg [7:0] out8131;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8131 = in0;
    end

    reg [7:0] out8132;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8132 = in0;
    end

    reg [7:0] out8133;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8133 = in0;
    end

    reg [7:0] out8134;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8134 = in0;
    end

    reg [7:0] out8135;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8135 = in0;
    end

    reg [7:0] out8136;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8136 = in0;
    end

    reg [7:0] out8137;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8137 = in0;
    end

    reg [7:0] out8138;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8138 = in0;
    end

    reg [7:0] out8139;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8139 = in0;
    end

    reg [7:0] out8140;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8140 = in0;
    end

    reg [7:0] out8141;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8141 = in0;
    end

    reg [7:0] out8142;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8142 = in0;
    end

    reg [7:0] out8143;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8143 = in0;
    end

    reg [7:0] out8144;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8144 = in0;
    end

    reg [7:0] out8145;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8145 = in0;
    end

    reg [7:0] out8146;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8146 = in0;
    end

    reg [7:0] out8147;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8147 = in0;
    end

    reg [7:0] out8148;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8148 = in0;
    end

    reg [7:0] out8149;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8149 = in0;
    end

    reg [7:0] out8150;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8150 = in0;
    end

    reg [7:0] out8151;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8151 = in0;
    end

    reg [7:0] out8152;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8152 = in0;
    end

    reg [7:0] out8153;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8153 = in0;
    end

    reg [7:0] out8154;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8154 = in0;
    end

    reg [7:0] out8155;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8155 = in0;
    end

    reg [7:0] out8156;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8156 = in0;
    end

    reg [7:0] out8157;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8157 = in0;
    end

    reg [7:0] out8158;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8158 = in0;
    end

    reg [7:0] out8159;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8159 = in0;
    end

    reg [7:0] out8160;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8160 = in0;
    end

    reg [7:0] out8161;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8161 = in0;
    end

    reg [7:0] out8162;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8162 = in0;
    end

    reg [7:0] out8163;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8163 = in0;
    end

    reg [7:0] out8164;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8164 = in0;
    end

    reg [7:0] out8165;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8165 = in0;
    end

    reg [7:0] out8166;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8166 = in0;
    end

    reg [7:0] out8167;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8167 = in0;
    end

    reg [7:0] out8168;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8168 = in0;
    end

    reg [7:0] out8169;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8169 = in0;
    end

    reg [7:0] out8170;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8170 = in0;
    end

    reg [7:0] out8171;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8171 = in0;
    end

    reg [7:0] out8172;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8172 = in0;
    end

    reg [7:0] out8173;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8173 = in0;
    end

    reg [7:0] out8174;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8174 = in0;
    end

    reg [7:0] out8175;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8175 = in0;
    end

    reg [7:0] out8176;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8176 = in0;
    end

    reg [7:0] out8177;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8177 = in0;
    end

    reg [7:0] out8178;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8178 = in0;
    end

    reg [7:0] out8179;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8179 = in0;
    end

    reg [7:0] out8180;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8180 = in0;
    end

    reg [7:0] out8181;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8181 = in0;
    end

    reg [7:0] out8182;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8182 = in0;
    end

    reg [7:0] out8183;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8183 = in0;
    end

    reg [7:0] out8184;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8184 = in0;
    end

    reg [7:0] out8185;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8185 = in0;
    end

    reg [7:0] out8186;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8186 = in0;
    end

    reg [7:0] out8187;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8187 = in0;
    end

    reg [7:0] out8188;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8188 = in0;
    end

    reg [7:0] out8189;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8189 = in0;
    end

    reg [7:0] out8190;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8190 = in0;
    end

    reg [7:0] out8191;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8191 = in0;
    end

    reg [7:0] out8192;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8192 = in0;
    end

    reg [7:0] out8193;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8193 = in0;
    end

    reg [7:0] out8194;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8194 = in0;
    end

    reg [7:0] out8195;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8195 = in0;
    end

    reg [7:0] out8196;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8196 = in0;
    end

    reg [7:0] out8197;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8197 = in0;
    end

    reg [7:0] out8198;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8198 = in0;
    end

    reg [7:0] out8199;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8199 = in0;
    end

    reg [7:0] out8200;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8200 = in0;
    end

    reg [7:0] out8201;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8201 = in0;
    end

    reg [7:0] out8202;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8202 = in0;
    end

    reg [7:0] out8203;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8203 = in0;
    end

    reg [7:0] out8204;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8204 = in0;
    end

    reg [7:0] out8205;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8205 = in0;
    end

    reg [7:0] out8206;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8206 = in0;
    end

    reg [7:0] out8207;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8207 = in0;
    end

    reg [7:0] out8208;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8208 = in0;
    end

    reg [7:0] out8209;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8209 = in0;
    end

    reg [7:0] out8210;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8210 = in0;
    end

    reg [7:0] out8211;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8211 = in0;
    end

    reg [7:0] out8212;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8212 = in0;
    end

    reg [7:0] out8213;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8213 = in0;
    end

    reg [7:0] out8214;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8214 = in0;
    end

    reg [7:0] out8215;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8215 = in0;
    end

    reg [7:0] out8216;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8216 = in0;
    end

    reg [7:0] out8217;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8217 = in0;
    end

    reg [7:0] out8218;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8218 = in0;
    end

    reg [7:0] out8219;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8219 = in0;
    end

    reg [7:0] out8220;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8220 = in0;
    end

    reg [7:0] out8221;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8221 = in0;
    end

    reg [7:0] out8222;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8222 = in0;
    end

    reg [7:0] out8223;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8223 = in0;
    end

    reg [7:0] out8224;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8224 = in0;
    end

    reg [7:0] out8225;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8225 = in0;
    end

    reg [7:0] out8226;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8226 = in0;
    end

    reg [7:0] out8227;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8227 = in0;
    end

    reg [7:0] out8228;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8228 = in0;
    end

    reg [7:0] out8229;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8229 = in0;
    end

    reg [7:0] out8230;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8230 = in0;
    end

    reg [7:0] out8231;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8231 = in0;
    end

    reg [7:0] out8232;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8232 = in0;
    end

    reg [7:0] out8233;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8233 = in0;
    end

    reg [7:0] out8234;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8234 = in0;
    end

    reg [7:0] out8235;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8235 = in0;
    end

    reg [7:0] out8236;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8236 = in0;
    end

    reg [7:0] out8237;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8237 = in0;
    end

    reg [7:0] out8238;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8238 = in0;
    end

    reg [7:0] out8239;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8239 = in0;
    end

    reg [7:0] out8240;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8240 = in0;
    end

    reg [7:0] out8241;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8241 = in0;
    end

    reg [7:0] out8242;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8242 = in0;
    end

    reg [7:0] out8243;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8243 = in0;
    end

    reg [7:0] out8244;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8244 = in0;
    end

    reg [7:0] out8245;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8245 = in0;
    end

    reg [7:0] out8246;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8246 = in0;
    end

    reg [7:0] out8247;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8247 = in0;
    end

    reg [7:0] out8248;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8248 = in0;
    end

    reg [7:0] out8249;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8249 = in0;
    end

    reg [7:0] out8250;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8250 = in0;
    end

    reg [7:0] out8251;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8251 = in0;
    end

    reg [7:0] out8252;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8252 = in0;
    end

    reg [7:0] out8253;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8253 = in0;
    end

    reg [7:0] out8254;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8254 = in0;
    end

    reg [7:0] out8255;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8255 = in0;
    end

    reg [7:0] out8256;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8256 = in0;
    end

    reg [7:0] out8257;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8257 = in0;
    end

    reg [7:0] out8258;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8258 = in0;
    end

    reg [7:0] out8259;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8259 = in0;
    end

    reg [7:0] out8260;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8260 = in0;
    end

    reg [7:0] out8261;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8261 = in0;
    end

    reg [7:0] out8262;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8262 = in0;
    end

    reg [7:0] out8263;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8263 = in0;
    end

    reg [7:0] out8264;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8264 = in0;
    end

    reg [7:0] out8265;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8265 = in0;
    end

    reg [7:0] out8266;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8266 = in0;
    end

    reg [7:0] out8267;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8267 = in0;
    end

    reg [7:0] out8268;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8268 = in0;
    end

    reg [7:0] out8269;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8269 = in0;
    end

    reg [7:0] out8270;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8270 = in0;
    end

    reg [7:0] out8271;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8271 = in0;
    end

    reg [7:0] out8272;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8272 = in0;
    end

    reg [7:0] out8273;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8273 = in0;
    end

    reg [7:0] out8274;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8274 = in0;
    end

    reg [7:0] out8275;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8275 = in0;
    end

    reg [7:0] out8276;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8276 = in0;
    end

    reg [7:0] out8277;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8277 = in0;
    end

    reg [7:0] out8278;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8278 = in0;
    end

    reg [7:0] out8279;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8279 = in0;
    end

    reg [7:0] out8280;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8280 = in0;
    end

    reg [7:0] out8281;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8281 = in0;
    end

    reg [7:0] out8282;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8282 = in0;
    end

    reg [7:0] out8283;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8283 = in0;
    end

    reg [7:0] out8284;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8284 = in0;
    end

    reg [7:0] out8285;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8285 = in0;
    end

    reg [7:0] out8286;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8286 = in0;
    end

    reg [7:0] out8287;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8287 = in0;
    end

    reg [7:0] out8288;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8288 = in0;
    end

    reg [7:0] out8289;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8289 = in0;
    end

    reg [7:0] out8290;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8290 = in0;
    end

    reg [7:0] out8291;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8291 = in0;
    end

    reg [7:0] out8292;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8292 = in0;
    end

    reg [7:0] out8293;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8293 = in0;
    end

    reg [7:0] out8294;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8294 = in0;
    end

    reg [7:0] out8295;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8295 = in0;
    end

    reg [7:0] out8296;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8296 = in0;
    end

    reg [7:0] out8297;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8297 = in0;
    end

    reg [7:0] out8298;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8298 = in0;
    end

    reg [7:0] out8299;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8299 = in0;
    end

    reg [7:0] out8300;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8300 = in0;
    end

    reg [7:0] out8301;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8301 = in0;
    end

    reg [7:0] out8302;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8302 = in0;
    end

    reg [7:0] out8303;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8303 = in0;
    end

    reg [7:0] out8304;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8304 = in0;
    end

    reg [7:0] out8305;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8305 = in0;
    end

    reg [7:0] out8306;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8306 = in0;
    end

    reg [7:0] out8307;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8307 = in0;
    end

    reg [7:0] out8308;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8308 = in0;
    end

    reg [7:0] out8309;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8309 = in0;
    end

    reg [7:0] out8310;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8310 = in0;
    end

    reg [7:0] out8311;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8311 = in0;
    end

    reg [7:0] out8312;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8312 = in0;
    end

    reg [7:0] out8313;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8313 = in0;
    end

    reg [7:0] out8314;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8314 = in0;
    end

    reg [7:0] out8315;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8315 = in0;
    end

    reg [7:0] out8316;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8316 = in0;
    end

    reg [7:0] out8317;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8317 = in0;
    end

    reg [7:0] out8318;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8318 = in0;
    end

    reg [7:0] out8319;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8319 = in0;
    end

    reg [7:0] out8320;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8320 = in0;
    end

    reg [7:0] out8321;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8321 = in0;
    end

    reg [7:0] out8322;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8322 = in0;
    end

    reg [7:0] out8323;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8323 = in0;
    end

    reg [7:0] out8324;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8324 = in0;
    end

    reg [7:0] out8325;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8325 = in0;
    end

    reg [7:0] out8326;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8326 = in0;
    end

    reg [7:0] out8327;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8327 = in0;
    end

    reg [7:0] out8328;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8328 = in0;
    end

    reg [7:0] out8329;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8329 = in0;
    end

    reg [7:0] out8330;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8330 = in0;
    end

    reg [7:0] out8331;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8331 = in0;
    end

    reg [7:0] out8332;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8332 = in0;
    end

    reg [7:0] out8333;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8333 = in0;
    end

    reg [7:0] out8334;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8334 = in0;
    end

    reg [7:0] out8335;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8335 = in0;
    end

    reg [7:0] out8336;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8336 = in0;
    end

    reg [7:0] out8337;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8337 = in0;
    end

    reg [7:0] out8338;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8338 = in0;
    end

    reg [7:0] out8339;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8339 = in0;
    end

    reg [7:0] out8340;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8340 = in0;
    end

    reg [7:0] out8341;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8341 = in0;
    end

    reg [7:0] out8342;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8342 = in0;
    end

    reg [7:0] out8343;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8343 = in0;
    end

    reg [7:0] out8344;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8344 = in0;
    end

    reg [7:0] out8345;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8345 = in0;
    end

    reg [7:0] out8346;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8346 = in0;
    end

    reg [7:0] out8347;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8347 = in0;
    end

    reg [7:0] out8348;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8348 = in0;
    end

    reg [7:0] out8349;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8349 = in0;
    end

    reg [7:0] out8350;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8350 = in0;
    end

    reg [7:0] out8351;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8351 = in0;
    end

    reg [7:0] out8352;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8352 = in0;
    end

    reg [7:0] out8353;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8353 = in0;
    end

    reg [7:0] out8354;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8354 = in0;
    end

    reg [7:0] out8355;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8355 = in0;
    end

    reg [7:0] out8356;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8356 = in0;
    end

    reg [7:0] out8357;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8357 = in0;
    end

    reg [7:0] out8358;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8358 = in0;
    end

    reg [7:0] out8359;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8359 = in0;
    end

    reg [7:0] out8360;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8360 = in0;
    end

    reg [7:0] out8361;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8361 = in0;
    end

    reg [7:0] out8362;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8362 = in0;
    end

    reg [7:0] out8363;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8363 = in0;
    end

    reg [7:0] out8364;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8364 = in0;
    end

    reg [7:0] out8365;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8365 = in0;
    end

    reg [7:0] out8366;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8366 = in0;
    end

    reg [7:0] out8367;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8367 = in0;
    end

    reg [7:0] out8368;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8368 = in0;
    end

    reg [7:0] out8369;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8369 = in0;
    end

    reg [7:0] out8370;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8370 = in0;
    end

    reg [7:0] out8371;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8371 = in0;
    end

    reg [7:0] out8372;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8372 = in0;
    end

    reg [7:0] out8373;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8373 = in0;
    end

    reg [7:0] out8374;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8374 = in0;
    end

    reg [7:0] out8375;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8375 = in0;
    end

    reg [7:0] out8376;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8376 = in0;
    end

    reg [7:0] out8377;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8377 = in0;
    end

    reg [7:0] out8378;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8378 = in0;
    end

    reg [7:0] out8379;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8379 = in0;
    end

    reg [7:0] out8380;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8380 = in0;
    end

    reg [7:0] out8381;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8381 = in0;
    end

    reg [7:0] out8382;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8382 = in0;
    end

    reg [7:0] out8383;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8383 = in0;
    end

    reg [7:0] out8384;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8384 = in0;
    end

    reg [7:0] out8385;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8385 = in0;
    end

    reg [7:0] out8386;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8386 = in0;
    end

    reg [7:0] out8387;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8387 = in0;
    end

    reg [7:0] out8388;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8388 = in0;
    end

    reg [7:0] out8389;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8389 = in0;
    end

    reg [7:0] out8390;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8390 = in0;
    end

    reg [7:0] out8391;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8391 = in0;
    end

    reg [7:0] out8392;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8392 = in0;
    end

    reg [7:0] out8393;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8393 = in0;
    end

    reg [7:0] out8394;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8394 = in0;
    end

    reg [7:0] out8395;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8395 = in0;
    end

    reg [7:0] out8396;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8396 = in0;
    end

    reg [7:0] out8397;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8397 = in0;
    end

    reg [7:0] out8398;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8398 = in0;
    end

    reg [7:0] out8399;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8399 = in0;
    end

    reg [7:0] out8400;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8400 = in0;
    end

    reg [7:0] out8401;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8401 = in0;
    end

    reg [7:0] out8402;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8402 = in0;
    end

    reg [7:0] out8403;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8403 = in0;
    end

    reg [7:0] out8404;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8404 = in0;
    end

    reg [7:0] out8405;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8405 = in0;
    end

    reg [7:0] out8406;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8406 = in0;
    end

    reg [7:0] out8407;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8407 = in0;
    end

    reg [7:0] out8408;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8408 = in0;
    end

    reg [7:0] out8409;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8409 = in0;
    end

    reg [7:0] out8410;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8410 = in0;
    end

    reg [7:0] out8411;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8411 = in0;
    end

    reg [7:0] out8412;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8412 = in0;
    end

    reg [7:0] out8413;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8413 = in0;
    end

    reg [7:0] out8414;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8414 = in0;
    end

    reg [7:0] out8415;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8415 = in0;
    end

    reg [7:0] out8416;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8416 = in0;
    end

    reg [7:0] out8417;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8417 = in0;
    end

    reg [7:0] out8418;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8418 = in0;
    end

    reg [7:0] out8419;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8419 = in0;
    end

    reg [7:0] out8420;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8420 = in0;
    end

    reg [7:0] out8421;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8421 = in0;
    end

    reg [7:0] out8422;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8422 = in0;
    end

    reg [7:0] out8423;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8423 = in0;
    end

    reg [7:0] out8424;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8424 = in0;
    end

    reg [7:0] out8425;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8425 = in0;
    end

    reg [7:0] out8426;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8426 = in0;
    end

    reg [7:0] out8427;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8427 = in0;
    end

    reg [7:0] out8428;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8428 = in0;
    end

    reg [7:0] out8429;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8429 = in0;
    end

    reg [7:0] out8430;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8430 = in0;
    end

    reg [7:0] out8431;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8431 = in0;
    end

    reg [7:0] out8432;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8432 = in0;
    end

    reg [7:0] out8433;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8433 = in0;
    end

    reg [7:0] out8434;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8434 = in0;
    end

    reg [7:0] out8435;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8435 = in0;
    end

    reg [7:0] out8436;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8436 = in0;
    end

    reg [7:0] out8437;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8437 = in0;
    end

    reg [7:0] out8438;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8438 = in0;
    end

    reg [7:0] out8439;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8439 = in0;
    end

    reg [7:0] out8440;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8440 = in0;
    end

    reg [7:0] out8441;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8441 = in0;
    end

    reg [7:0] out8442;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8442 = in0;
    end

    reg [7:0] out8443;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8443 = in0;
    end

    reg [7:0] out8444;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8444 = in0;
    end

    reg [7:0] out8445;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8445 = in0;
    end

    reg [7:0] out8446;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8446 = in0;
    end

    reg [7:0] out8447;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8447 = in0;
    end

    reg [7:0] out8448;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8448 = in0;
    end

    reg [7:0] out8449;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8449 = in0;
    end

    reg [7:0] out8450;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8450 = in0;
    end

    reg [7:0] out8451;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8451 = in0;
    end

    reg [7:0] out8452;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8452 = in0;
    end

    reg [7:0] out8453;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8453 = in0;
    end

    reg [7:0] out8454;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8454 = in0;
    end

    reg [7:0] out8455;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8455 = in0;
    end

    reg [7:0] out8456;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8456 = in0;
    end

    reg [7:0] out8457;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8457 = in0;
    end

    reg [7:0] out8458;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8458 = in0;
    end

    reg [7:0] out8459;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8459 = in0;
    end

    reg [7:0] out8460;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8460 = in0;
    end

    reg [7:0] out8461;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8461 = in0;
    end

    reg [7:0] out8462;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8462 = in0;
    end

    reg [7:0] out8463;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8463 = in0;
    end

    reg [7:0] out8464;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8464 = in0;
    end

    reg [7:0] out8465;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8465 = in0;
    end

    reg [7:0] out8466;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8466 = in0;
    end

    reg [7:0] out8467;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8467 = in0;
    end

    reg [7:0] out8468;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8468 = in0;
    end

    reg [7:0] out8469;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8469 = in0;
    end

    reg [7:0] out8470;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8470 = in0;
    end

    reg [7:0] out8471;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8471 = in0;
    end

    reg [7:0] out8472;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8472 = in0;
    end

    reg [7:0] out8473;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8473 = in0;
    end

    reg [7:0] out8474;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8474 = in0;
    end

    reg [7:0] out8475;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8475 = in0;
    end

    reg [7:0] out8476;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8476 = in0;
    end

    reg [7:0] out8477;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8477 = in0;
    end

    reg [7:0] out8478;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8478 = in0;
    end

    reg [7:0] out8479;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8479 = in0;
    end

    reg [7:0] out8480;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8480 = in0;
    end

    reg [7:0] out8481;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8481 = in0;
    end

    reg [7:0] out8482;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8482 = in0;
    end

    reg [7:0] out8483;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8483 = in0;
    end

    reg [7:0] out8484;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8484 = in0;
    end

    reg [7:0] out8485;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8485 = in0;
    end

    reg [7:0] out8486;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8486 = in0;
    end

    reg [7:0] out8487;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8487 = in0;
    end

    reg [7:0] out8488;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8488 = in0;
    end

    reg [7:0] out8489;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8489 = in0;
    end

    reg [7:0] out8490;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8490 = in0;
    end

    reg [7:0] out8491;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8491 = in0;
    end

    reg [7:0] out8492;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8492 = in0;
    end

    reg [7:0] out8493;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8493 = in0;
    end

    reg [7:0] out8494;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8494 = in0;
    end

    reg [7:0] out8495;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8495 = in0;
    end

    reg [7:0] out8496;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8496 = in0;
    end

    reg [7:0] out8497;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8497 = in0;
    end

    reg [7:0] out8498;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8498 = in0;
    end

    reg [7:0] out8499;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8499 = in0;
    end

    reg [7:0] out8500;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8500 = in0;
    end

    reg [7:0] out8501;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8501 = in0;
    end

    reg [7:0] out8502;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8502 = in0;
    end

    reg [7:0] out8503;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8503 = in0;
    end

    reg [7:0] out8504;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8504 = in0;
    end

    reg [7:0] out8505;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8505 = in0;
    end

    reg [7:0] out8506;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8506 = in0;
    end

    reg [7:0] out8507;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8507 = in0;
    end

    reg [7:0] out8508;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8508 = in0;
    end

    reg [7:0] out8509;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8509 = in0;
    end

    reg [7:0] out8510;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8510 = in0;
    end

    reg [7:0] out8511;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8511 = in0;
    end

    reg [7:0] out8512;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8512 = in0;
    end

    reg [7:0] out8513;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8513 = in0;
    end

    reg [7:0] out8514;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8514 = in0;
    end

    reg [7:0] out8515;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8515 = in0;
    end

    reg [7:0] out8516;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8516 = in0;
    end

    reg [7:0] out8517;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8517 = in0;
    end

    reg [7:0] out8518;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8518 = in0;
    end

    reg [7:0] out8519;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8519 = in0;
    end

    reg [7:0] out8520;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8520 = in0;
    end

    reg [7:0] out8521;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8521 = in0;
    end

    reg [7:0] out8522;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8522 = in0;
    end

    reg [7:0] out8523;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8523 = in0;
    end

    reg [7:0] out8524;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8524 = in0;
    end

    reg [7:0] out8525;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8525 = in0;
    end

    reg [7:0] out8526;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8526 = in0;
    end

    reg [7:0] out8527;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8527 = in0;
    end

    reg [7:0] out8528;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8528 = in0;
    end

    reg [7:0] out8529;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8529 = in0;
    end

    reg [7:0] out8530;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8530 = in0;
    end

    reg [7:0] out8531;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8531 = in0;
    end

    reg [7:0] out8532;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8532 = in0;
    end

    reg [7:0] out8533;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8533 = in0;
    end

    reg [7:0] out8534;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8534 = in0;
    end

    reg [7:0] out8535;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8535 = in0;
    end

    reg [7:0] out8536;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8536 = in0;
    end

    reg [7:0] out8537;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8537 = in0;
    end

    reg [7:0] out8538;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8538 = in0;
    end

    reg [7:0] out8539;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8539 = in0;
    end

    reg [7:0] out8540;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8540 = in0;
    end

    reg [7:0] out8541;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8541 = in0;
    end

    reg [7:0] out8542;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8542 = in0;
    end

    reg [7:0] out8543;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8543 = in0;
    end

    reg [7:0] out8544;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8544 = in0;
    end

    reg [7:0] out8545;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8545 = in0;
    end

    reg [7:0] out8546;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8546 = in0;
    end

    reg [7:0] out8547;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8547 = in0;
    end

    reg [7:0] out8548;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8548 = in0;
    end

    reg [7:0] out8549;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8549 = in0;
    end

    reg [7:0] out8550;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8550 = in0;
    end

    reg [7:0] out8551;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8551 = in0;
    end

    reg [7:0] out8552;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8552 = in0;
    end

    reg [7:0] out8553;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8553 = in0;
    end

    reg [7:0] out8554;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8554 = in0;
    end

    reg [7:0] out8555;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8555 = in0;
    end

    reg [7:0] out8556;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8556 = in0;
    end

    reg [7:0] out8557;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8557 = in0;
    end

    reg [7:0] out8558;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8558 = in0;
    end

    reg [7:0] out8559;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8559 = in0;
    end

    reg [7:0] out8560;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8560 = in0;
    end

    reg [7:0] out8561;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8561 = in0;
    end

    reg [7:0] out8562;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8562 = in0;
    end

    reg [7:0] out8563;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8563 = in0;
    end

    reg [7:0] out8564;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8564 = in0;
    end

    reg [7:0] out8565;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8565 = in0;
    end

    reg [7:0] out8566;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8566 = in0;
    end

    reg [7:0] out8567;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8567 = in0;
    end

    reg [7:0] out8568;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8568 = in0;
    end

    reg [7:0] out8569;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8569 = in0;
    end

    reg [7:0] out8570;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8570 = in0;
    end

    reg [7:0] out8571;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8571 = in0;
    end

    reg [7:0] out8572;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8572 = in0;
    end

    reg [7:0] out8573;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8573 = in0;
    end

    reg [7:0] out8574;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8574 = in0;
    end

    reg [7:0] out8575;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8575 = in0;
    end

    reg [7:0] out8576;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8576 = in0;
    end

    reg [7:0] out8577;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8577 = in0;
    end

    reg [7:0] out8578;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8578 = in0;
    end

    reg [7:0] out8579;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8579 = in0;
    end

    reg [7:0] out8580;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8580 = in0;
    end

    reg [7:0] out8581;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8581 = in0;
    end

    reg [7:0] out8582;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8582 = in0;
    end

    reg [7:0] out8583;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8583 = in0;
    end

    reg [7:0] out8584;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8584 = in0;
    end

    reg [7:0] out8585;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8585 = in0;
    end

    reg [7:0] out8586;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8586 = in0;
    end

    reg [7:0] out8587;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8587 = in0;
    end

    reg [7:0] out8588;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8588 = in0;
    end

    reg [7:0] out8589;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8589 = in0;
    end

    reg [7:0] out8590;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8590 = in0;
    end

    reg [7:0] out8591;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8591 = in0;
    end

    reg [7:0] out8592;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8592 = in0;
    end

    reg [7:0] out8593;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8593 = in0;
    end

    reg [7:0] out8594;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8594 = in0;
    end

    reg [7:0] out8595;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8595 = in0;
    end

    reg [7:0] out8596;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8596 = in0;
    end

    reg [7:0] out8597;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8597 = in0;
    end

    reg [7:0] out8598;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8598 = in0;
    end

    reg [7:0] out8599;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8599 = in0;
    end

    reg [7:0] out8600;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8600 = in0;
    end

    reg [7:0] out8601;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8601 = in0;
    end

    reg [7:0] out8602;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8602 = in0;
    end

    reg [7:0] out8603;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8603 = in0;
    end

    reg [7:0] out8604;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8604 = in0;
    end

    reg [7:0] out8605;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8605 = in0;
    end

    reg [7:0] out8606;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8606 = in0;
    end

    reg [7:0] out8607;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8607 = in0;
    end

    reg [7:0] out8608;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8608 = in0;
    end

    reg [7:0] out8609;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8609 = in0;
    end

    reg [7:0] out8610;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8610 = in0;
    end

    reg [7:0] out8611;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8611 = in0;
    end

    reg [7:0] out8612;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8612 = in0;
    end

    reg [7:0] out8613;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8613 = in0;
    end

    reg [7:0] out8614;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8614 = in0;
    end

    reg [7:0] out8615;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8615 = in0;
    end

    reg [7:0] out8616;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8616 = in0;
    end

    reg [7:0] out8617;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8617 = in0;
    end

    reg [7:0] out8618;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8618 = in0;
    end

    reg [7:0] out8619;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8619 = in0;
    end

    reg [7:0] out8620;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8620 = in0;
    end

    reg [7:0] out8621;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8621 = in0;
    end

    reg [7:0] out8622;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8622 = in0;
    end

    reg [7:0] out8623;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8623 = in0;
    end

    reg [7:0] out8624;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8624 = in0;
    end

    reg [7:0] out8625;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8625 = in0;
    end

    reg [7:0] out8626;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8626 = in0;
    end

    reg [7:0] out8627;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8627 = in0;
    end

    reg [7:0] out8628;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8628 = in0;
    end

    reg [7:0] out8629;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8629 = in0;
    end

    reg [7:0] out8630;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8630 = in0;
    end

    reg [7:0] out8631;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8631 = in0;
    end

    reg [7:0] out8632;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8632 = in0;
    end

    reg [7:0] out8633;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8633 = in0;
    end

    reg [7:0] out8634;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8634 = in0;
    end

    reg [7:0] out8635;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8635 = in0;
    end

    reg [7:0] out8636;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8636 = in0;
    end

    reg [7:0] out8637;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8637 = in0;
    end

    reg [7:0] out8638;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8638 = in0;
    end

    reg [7:0] out8639;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8639 = in0;
    end

    reg [7:0] out8640;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8640 = in0;
    end

    reg [7:0] out8641;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8641 = in0;
    end

    reg [7:0] out8642;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8642 = in0;
    end

    reg [7:0] out8643;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8643 = in0;
    end

    reg [7:0] out8644;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8644 = in0;
    end

    reg [7:0] out8645;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8645 = in0;
    end

    reg [7:0] out8646;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8646 = in0;
    end

    reg [7:0] out8647;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8647 = in0;
    end

    reg [7:0] out8648;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8648 = in0;
    end

    reg [7:0] out8649;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8649 = in0;
    end

    reg [7:0] out8650;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8650 = in0;
    end

    reg [7:0] out8651;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8651 = in0;
    end

    reg [7:0] out8652;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8652 = in0;
    end

    reg [7:0] out8653;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8653 = in0;
    end

    reg [7:0] out8654;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8654 = in0;
    end

    reg [7:0] out8655;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8655 = in0;
    end

    reg [7:0] out8656;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8656 = in0;
    end

    reg [7:0] out8657;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8657 = in0;
    end

    reg [7:0] out8658;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8658 = in0;
    end

    reg [7:0] out8659;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8659 = in0;
    end

    reg [7:0] out8660;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8660 = in0;
    end

    reg [7:0] out8661;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8661 = in0;
    end

    reg [7:0] out8662;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8662 = in0;
    end

    reg [7:0] out8663;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8663 = in0;
    end

    reg [7:0] out8664;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8664 = in0;
    end

    reg [7:0] out8665;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8665 = in0;
    end

    reg [7:0] out8666;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8666 = in0;
    end

    reg [7:0] out8667;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8667 = in0;
    end

    reg [7:0] out8668;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8668 = in0;
    end

    reg [7:0] out8669;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8669 = in0;
    end

    reg [7:0] out8670;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8670 = in0;
    end

    reg [7:0] out8671;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8671 = in0;
    end

    reg [7:0] out8672;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8672 = in0;
    end

    reg [7:0] out8673;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8673 = in0;
    end

    reg [7:0] out8674;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8674 = in0;
    end

    reg [7:0] out8675;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8675 = in0;
    end

    reg [7:0] out8676;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8676 = in0;
    end

    reg [7:0] out8677;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8677 = in0;
    end

    reg [7:0] out8678;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8678 = in0;
    end

    reg [7:0] out8679;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8679 = in0;
    end

    reg [7:0] out8680;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8680 = in0;
    end

    reg [7:0] out8681;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8681 = in0;
    end

    reg [7:0] out8682;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8682 = in0;
    end

    reg [7:0] out8683;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8683 = in0;
    end

    reg [7:0] out8684;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8684 = in0;
    end

    reg [7:0] out8685;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8685 = in0;
    end

    reg [7:0] out8686;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8686 = in0;
    end

    reg [7:0] out8687;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8687 = in0;
    end

    reg [7:0] out8688;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8688 = in0;
    end

    reg [7:0] out8689;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8689 = in0;
    end

    reg [7:0] out8690;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8690 = in0;
    end

    reg [7:0] out8691;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8691 = in0;
    end

    reg [7:0] out8692;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8692 = in0;
    end

    reg [7:0] out8693;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8693 = in0;
    end

    reg [7:0] out8694;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8694 = in0;
    end

    reg [7:0] out8695;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8695 = in0;
    end

    reg [7:0] out8696;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8696 = in0;
    end

    reg [7:0] out8697;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8697 = in0;
    end

    reg [7:0] out8698;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8698 = in0;
    end

    reg [7:0] out8699;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8699 = in0;
    end

    reg [7:0] out8700;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8700 = in0;
    end

    reg [7:0] out8701;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8701 = in0;
    end

    reg [7:0] out8702;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8702 = in0;
    end

    reg [7:0] out8703;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8703 = in0;
    end

    reg [7:0] out8704;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8704 = in0;
    end

    reg [7:0] out8705;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8705 = in0;
    end

    reg [7:0] out8706;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8706 = in0;
    end

    reg [7:0] out8707;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8707 = in0;
    end

    reg [7:0] out8708;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8708 = in0;
    end

    reg [7:0] out8709;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8709 = in0;
    end

    reg [7:0] out8710;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8710 = in0;
    end

    reg [7:0] out8711;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8711 = in0;
    end

    reg [7:0] out8712;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8712 = in0;
    end

    reg [7:0] out8713;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8713 = in0;
    end

    reg [7:0] out8714;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8714 = in0;
    end

    reg [7:0] out8715;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8715 = in0;
    end

    reg [7:0] out8716;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8716 = in0;
    end

    reg [7:0] out8717;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8717 = in0;
    end

    reg [7:0] out8718;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8718 = in0;
    end

    reg [7:0] out8719;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8719 = in0;
    end

    reg [7:0] out8720;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8720 = in0;
    end

    reg [7:0] out8721;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8721 = in0;
    end

    reg [7:0] out8722;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8722 = in0;
    end

    reg [7:0] out8723;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8723 = in0;
    end

    reg [7:0] out8724;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8724 = in0;
    end

    reg [7:0] out8725;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8725 = in0;
    end

    reg [7:0] out8726;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8726 = in0;
    end

    reg [7:0] out8727;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8727 = in0;
    end

    reg [7:0] out8728;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8728 = in0;
    end

    reg [7:0] out8729;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8729 = in0;
    end

    reg [7:0] out8730;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8730 = in0;
    end

    reg [7:0] out8731;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8731 = in0;
    end

    reg [7:0] out8732;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8732 = in0;
    end

    reg [7:0] out8733;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8733 = in0;
    end

    reg [7:0] out8734;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8734 = in0;
    end

    reg [7:0] out8735;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8735 = in0;
    end

    reg [7:0] out8736;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8736 = in0;
    end

    reg [7:0] out8737;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8737 = in0;
    end

    reg [7:0] out8738;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8738 = in0;
    end

    reg [7:0] out8739;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8739 = in0;
    end

    reg [7:0] out8740;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8740 = in0;
    end

    reg [7:0] out8741;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8741 = in0;
    end

    reg [7:0] out8742;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8742 = in0;
    end

    reg [7:0] out8743;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8743 = in0;
    end

    reg [7:0] out8744;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8744 = in0;
    end

    reg [7:0] out8745;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8745 = in0;
    end

    reg [7:0] out8746;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8746 = in0;
    end

    reg [7:0] out8747;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8747 = in0;
    end

    reg [7:0] out8748;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8748 = in0;
    end

    reg [7:0] out8749;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8749 = in0;
    end

    reg [7:0] out8750;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8750 = in0;
    end

    reg [7:0] out8751;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8751 = in0;
    end

    reg [7:0] out8752;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8752 = in0;
    end

    reg [7:0] out8753;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8753 = in0;
    end

    reg [7:0] out8754;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8754 = in0;
    end

    reg [7:0] out8755;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8755 = in0;
    end

    reg [7:0] out8756;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8756 = in0;
    end

    reg [7:0] out8757;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8757 = in0;
    end

    reg [7:0] out8758;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8758 = in0;
    end

    reg [7:0] out8759;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8759 = in0;
    end

    reg [7:0] out8760;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8760 = in0;
    end

    reg [7:0] out8761;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8761 = in0;
    end

    reg [7:0] out8762;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8762 = in0;
    end

    reg [7:0] out8763;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8763 = in0;
    end

    reg [7:0] out8764;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8764 = in0;
    end

    reg [7:0] out8765;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8765 = in0;
    end

    reg [7:0] out8766;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8766 = in0;
    end

    reg [7:0] out8767;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8767 = in0;
    end

    reg [7:0] out8768;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8768 = in0;
    end

    reg [7:0] out8769;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8769 = in0;
    end

    reg [7:0] out8770;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8770 = in0;
    end

    reg [7:0] out8771;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8771 = in0;
    end

    reg [7:0] out8772;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8772 = in0;
    end

    reg [7:0] out8773;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8773 = in0;
    end

    reg [7:0] out8774;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8774 = in0;
    end

    reg [7:0] out8775;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8775 = in0;
    end

    reg [7:0] out8776;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8776 = in0;
    end

    reg [7:0] out8777;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8777 = in0;
    end

    reg [7:0] out8778;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8778 = in0;
    end

    reg [7:0] out8779;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8779 = in0;
    end

    reg [7:0] out8780;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8780 = in0;
    end

    reg [7:0] out8781;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8781 = in0;
    end

    reg [7:0] out8782;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8782 = in0;
    end

    reg [7:0] out8783;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8783 = in0;
    end

    reg [7:0] out8784;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8784 = in0;
    end

    reg [7:0] out8785;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8785 = in0;
    end

    reg [7:0] out8786;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8786 = in0;
    end

    reg [7:0] out8787;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8787 = in0;
    end

    reg [7:0] out8788;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8788 = in0;
    end

    reg [7:0] out8789;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8789 = in0;
    end

    reg [7:0] out8790;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8790 = in0;
    end

    reg [7:0] out8791;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8791 = in0;
    end

    reg [7:0] out8792;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8792 = in0;
    end

    reg [7:0] out8793;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8793 = in0;
    end

    reg [7:0] out8794;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8794 = in0;
    end

    reg [7:0] out8795;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8795 = in0;
    end

    reg [7:0] out8796;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8796 = in0;
    end

    reg [7:0] out8797;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8797 = in0;
    end

    reg [7:0] out8798;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8798 = in0;
    end

    reg [7:0] out8799;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8799 = in0;
    end

    reg [7:0] out8800;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8800 = in0;
    end

    reg [7:0] out8801;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8801 = in0;
    end

    reg [7:0] out8802;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8802 = in0;
    end

    reg [7:0] out8803;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8803 = in0;
    end

    reg [7:0] out8804;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8804 = in0;
    end

    reg [7:0] out8805;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8805 = in0;
    end

    reg [7:0] out8806;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8806 = in0;
    end

    reg [7:0] out8807;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8807 = in0;
    end

    reg [7:0] out8808;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8808 = in0;
    end

    reg [7:0] out8809;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8809 = in0;
    end

    reg [7:0] out8810;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8810 = in0;
    end

    reg [7:0] out8811;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8811 = in0;
    end

    reg [7:0] out8812;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8812 = in0;
    end

    reg [7:0] out8813;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8813 = in0;
    end

    reg [7:0] out8814;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8814 = in0;
    end

    reg [7:0] out8815;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8815 = in0;
    end

    reg [7:0] out8816;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8816 = in0;
    end

    reg [7:0] out8817;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8817 = in0;
    end

    reg [7:0] out8818;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8818 = in0;
    end

    reg [7:0] out8819;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8819 = in0;
    end

    reg [7:0] out8820;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8820 = in0;
    end

    reg [7:0] out8821;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8821 = in0;
    end

    reg [7:0] out8822;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8822 = in0;
    end

    reg [7:0] out8823;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8823 = in0;
    end

    reg [7:0] out8824;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8824 = in0;
    end

    reg [7:0] out8825;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8825 = in0;
    end

    reg [7:0] out8826;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8826 = in0;
    end

    reg [7:0] out8827;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8827 = in0;
    end

    reg [7:0] out8828;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8828 = in0;
    end

    reg [7:0] out8829;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8829 = in0;
    end

    reg [7:0] out8830;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8830 = in0;
    end

    reg [7:0] out8831;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8831 = in0;
    end

    reg [7:0] out8832;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8832 = in0;
    end

    reg [7:0] out8833;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8833 = in0;
    end

    reg [7:0] out8834;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8834 = in0;
    end

    reg [7:0] out8835;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8835 = in0;
    end

    reg [7:0] out8836;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8836 = in0;
    end

    reg [7:0] out8837;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8837 = in0;
    end

    reg [7:0] out8838;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8838 = in0;
    end

    reg [7:0] out8839;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8839 = in0;
    end

    reg [7:0] out8840;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8840 = in0;
    end

    reg [7:0] out8841;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8841 = in0;
    end

    reg [7:0] out8842;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8842 = in0;
    end

    reg [7:0] out8843;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8843 = in0;
    end

    reg [7:0] out8844;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8844 = in0;
    end

    reg [7:0] out8845;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8845 = in0;
    end

    reg [7:0] out8846;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8846 = in0;
    end

    reg [7:0] out8847;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8847 = in0;
    end

    reg [7:0] out8848;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8848 = in0;
    end

    reg [7:0] out8849;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8849 = in0;
    end

    reg [7:0] out8850;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8850 = in0;
    end

    reg [7:0] out8851;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8851 = in0;
    end

    reg [7:0] out8852;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8852 = in0;
    end

    reg [7:0] out8853;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8853 = in0;
    end

    reg [7:0] out8854;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8854 = in0;
    end

    reg [7:0] out8855;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8855 = in0;
    end

    reg [7:0] out8856;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8856 = in0;
    end

    reg [7:0] out8857;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8857 = in0;
    end

    reg [7:0] out8858;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8858 = in0;
    end

    reg [7:0] out8859;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8859 = in0;
    end

    reg [7:0] out8860;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8860 = in0;
    end

    reg [7:0] out8861;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8861 = in0;
    end

    reg [7:0] out8862;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8862 = in0;
    end

    reg [7:0] out8863;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8863 = in0;
    end

    reg [7:0] out8864;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8864 = in0;
    end

    reg [7:0] out8865;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8865 = in0;
    end

    reg [7:0] out8866;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8866 = in0;
    end

    reg [7:0] out8867;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8867 = in0;
    end

    reg [7:0] out8868;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8868 = in0;
    end

    reg [7:0] out8869;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8869 = in0;
    end

    reg [7:0] out8870;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8870 = in0;
    end

    reg [7:0] out8871;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8871 = in0;
    end

    reg [7:0] out8872;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8872 = in0;
    end

    reg [7:0] out8873;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8873 = in0;
    end

    reg [7:0] out8874;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8874 = in0;
    end

    reg [7:0] out8875;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8875 = in0;
    end

    reg [7:0] out8876;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8876 = in0;
    end

    reg [7:0] out8877;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8877 = in0;
    end

    reg [7:0] out8878;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8878 = in0;
    end

    reg [7:0] out8879;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8879 = in0;
    end

    reg [7:0] out8880;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8880 = in0;
    end

    reg [7:0] out8881;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8881 = in0;
    end

    reg [7:0] out8882;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8882 = in0;
    end

    reg [7:0] out8883;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8883 = in0;
    end

    reg [7:0] out8884;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8884 = in0;
    end

    reg [7:0] out8885;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8885 = in0;
    end

    reg [7:0] out8886;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8886 = in0;
    end

    reg [7:0] out8887;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8887 = in0;
    end

    reg [7:0] out8888;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8888 = in0;
    end

    reg [7:0] out8889;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8889 = in0;
    end

    reg [7:0] out8890;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8890 = in0;
    end

    reg [7:0] out8891;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8891 = in0;
    end

    reg [7:0] out8892;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8892 = in0;
    end

    reg [7:0] out8893;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8893 = in0;
    end

    reg [7:0] out8894;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8894 = in0;
    end

    reg [7:0] out8895;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8895 = in0;
    end

    reg [7:0] out8896;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8896 = in0;
    end

    reg [7:0] out8897;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8897 = in0;
    end

    reg [7:0] out8898;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8898 = in0;
    end

    reg [7:0] out8899;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8899 = in0;
    end

    reg [7:0] out8900;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8900 = in0;
    end

    reg [7:0] out8901;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8901 = in0;
    end

    reg [7:0] out8902;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8902 = in0;
    end

    reg [7:0] out8903;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8903 = in0;
    end

    reg [7:0] out8904;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8904 = in0;
    end

    reg [7:0] out8905;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8905 = in0;
    end

    reg [7:0] out8906;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8906 = in0;
    end

    reg [7:0] out8907;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8907 = in0;
    end

    reg [7:0] out8908;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8908 = in0;
    end

    reg [7:0] out8909;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8909 = in0;
    end

    reg [7:0] out8910;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8910 = in0;
    end

    reg [7:0] out8911;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8911 = in0;
    end

    reg [7:0] out8912;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8912 = in0;
    end

    reg [7:0] out8913;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8913 = in0;
    end

    reg [7:0] out8914;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8914 = in0;
    end

    reg [7:0] out8915;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8915 = in0;
    end

    reg [7:0] out8916;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8916 = in0;
    end

    reg [7:0] out8917;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8917 = in0;
    end

    reg [7:0] out8918;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8918 = in0;
    end

    reg [7:0] out8919;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8919 = in0;
    end

    reg [7:0] out8920;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8920 = in0;
    end

    reg [7:0] out8921;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8921 = in0;
    end

    reg [7:0] out8922;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8922 = in0;
    end

    reg [7:0] out8923;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8923 = in0;
    end

    reg [7:0] out8924;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8924 = in0;
    end

    reg [7:0] out8925;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8925 = in0;
    end

    reg [7:0] out8926;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8926 = in0;
    end

    reg [7:0] out8927;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8927 = in0;
    end

    reg [7:0] out8928;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8928 = in0;
    end

    reg [7:0] out8929;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8929 = in0;
    end

    reg [7:0] out8930;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8930 = in0;
    end

    reg [7:0] out8931;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8931 = in0;
    end

    reg [7:0] out8932;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8932 = in0;
    end

    reg [7:0] out8933;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8933 = in0;
    end

    reg [7:0] out8934;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8934 = in0;
    end

    reg [7:0] out8935;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8935 = in0;
    end

    reg [7:0] out8936;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8936 = in0;
    end

    reg [7:0] out8937;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8937 = in0;
    end

    reg [7:0] out8938;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8938 = in0;
    end

    reg [7:0] out8939;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8939 = in0;
    end

    reg [7:0] out8940;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8940 = in0;
    end

    reg [7:0] out8941;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8941 = in0;
    end

    reg [7:0] out8942;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8942 = in0;
    end

    reg [7:0] out8943;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8943 = in0;
    end

    reg [7:0] out8944;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8944 = in0;
    end

    reg [7:0] out8945;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8945 = in0;
    end

    reg [7:0] out8946;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8946 = in0;
    end

    reg [7:0] out8947;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8947 = in0;
    end

    reg [7:0] out8948;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8948 = in0;
    end

    reg [7:0] out8949;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8949 = in0;
    end

    reg [7:0] out8950;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8950 = in0;
    end

    reg [7:0] out8951;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8951 = in0;
    end

    reg [7:0] out8952;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8952 = in0;
    end

    reg [7:0] out8953;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8953 = in0;
    end

    reg [7:0] out8954;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8954 = in0;
    end

    reg [7:0] out8955;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8955 = in0;
    end

    reg [7:0] out8956;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8956 = in0;
    end

    reg [7:0] out8957;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8957 = in0;
    end

    reg [7:0] out8958;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8958 = in0;
    end

    reg [7:0] out8959;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8959 = in0;
    end

    reg [7:0] out8960;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8960 = in0;
    end

    reg [7:0] out8961;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8961 = in0;
    end

    reg [7:0] out8962;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8962 = in0;
    end

    reg [7:0] out8963;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8963 = in0;
    end

    reg [7:0] out8964;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8964 = in0;
    end

    reg [7:0] out8965;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8965 = in0;
    end

    reg [7:0] out8966;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8966 = in0;
    end

    reg [7:0] out8967;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8967 = in0;
    end

    reg [7:0] out8968;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8968 = in0;
    end

    reg [7:0] out8969;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8969 = in0;
    end

    reg [7:0] out8970;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8970 = in0;
    end

    reg [7:0] out8971;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8971 = in0;
    end

    reg [7:0] out8972;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8972 = in0;
    end

    reg [7:0] out8973;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8973 = in0;
    end

    reg [7:0] out8974;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8974 = in0;
    end

    reg [7:0] out8975;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8975 = in0;
    end

    reg [7:0] out8976;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8976 = in0;
    end

    reg [7:0] out8977;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8977 = in0;
    end

    reg [7:0] out8978;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8978 = in0;
    end

    reg [7:0] out8979;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8979 = in0;
    end

    reg [7:0] out8980;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8980 = in0;
    end

    reg [7:0] out8981;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8981 = in0;
    end

    reg [7:0] out8982;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8982 = in0;
    end

    reg [7:0] out8983;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8983 = in0;
    end

    reg [7:0] out8984;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8984 = in0;
    end

    reg [7:0] out8985;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8985 = in0;
    end

    reg [7:0] out8986;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8986 = in0;
    end

    reg [7:0] out8987;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8987 = in0;
    end

    reg [7:0] out8988;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8988 = in0;
    end

    reg [7:0] out8989;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8989 = in0;
    end

    reg [7:0] out8990;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8990 = in0;
    end

    reg [7:0] out8991;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8991 = in0;
    end

    reg [7:0] out8992;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8992 = in0;
    end

    reg [7:0] out8993;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8993 = in0;
    end

    reg [7:0] out8994;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8994 = in0;
    end

    reg [7:0] out8995;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8995 = in0;
    end

    reg [7:0] out8996;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8996 = in0;
    end

    reg [7:0] out8997;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8997 = in0;
    end

    reg [7:0] out8998;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8998 = in0;
    end

    reg [7:0] out8999;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out8999 = in0;
    end

    reg [7:0] out9000;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9000 = in0;
    end

    reg [7:0] out9001;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9001 = in0;
    end

    reg [7:0] out9002;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9002 = in0;
    end

    reg [7:0] out9003;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9003 = in0;
    end

    reg [7:0] out9004;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9004 = in0;
    end

    reg [7:0] out9005;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9005 = in0;
    end

    reg [7:0] out9006;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9006 = in0;
    end

    reg [7:0] out9007;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9007 = in0;
    end

    reg [7:0] out9008;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9008 = in0;
    end

    reg [7:0] out9009;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9009 = in0;
    end

    reg [7:0] out9010;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9010 = in0;
    end

    reg [7:0] out9011;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9011 = in0;
    end

    reg [7:0] out9012;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9012 = in0;
    end

    reg [7:0] out9013;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9013 = in0;
    end

    reg [7:0] out9014;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9014 = in0;
    end

    reg [7:0] out9015;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9015 = in0;
    end

    reg [7:0] out9016;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9016 = in0;
    end

    reg [7:0] out9017;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9017 = in0;
    end

    reg [7:0] out9018;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9018 = in0;
    end

    reg [7:0] out9019;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9019 = in0;
    end

    reg [7:0] out9020;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9020 = in0;
    end

    reg [7:0] out9021;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9021 = in0;
    end

    reg [7:0] out9022;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9022 = in0;
    end

    reg [7:0] out9023;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9023 = in0;
    end

    reg [7:0] out9024;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9024 = in0;
    end

    reg [7:0] out9025;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9025 = in0;
    end

    reg [7:0] out9026;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9026 = in0;
    end

    reg [7:0] out9027;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9027 = in0;
    end

    reg [7:0] out9028;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9028 = in0;
    end

    reg [7:0] out9029;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9029 = in0;
    end

    reg [7:0] out9030;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9030 = in0;
    end

    reg [7:0] out9031;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9031 = in0;
    end

    reg [7:0] out9032;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9032 = in0;
    end

    reg [7:0] out9033;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9033 = in0;
    end

    reg [7:0] out9034;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9034 = in0;
    end

    reg [7:0] out9035;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9035 = in0;
    end

    reg [7:0] out9036;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9036 = in0;
    end

    reg [7:0] out9037;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9037 = in0;
    end

    reg [7:0] out9038;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9038 = in0;
    end

    reg [7:0] out9039;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9039 = in0;
    end

    reg [7:0] out9040;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9040 = in0;
    end

    reg [7:0] out9041;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9041 = in0;
    end

    reg [7:0] out9042;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9042 = in0;
    end

    reg [7:0] out9043;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9043 = in0;
    end

    reg [7:0] out9044;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9044 = in0;
    end

    reg [7:0] out9045;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9045 = in0;
    end

    reg [7:0] out9046;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9046 = in0;
    end

    reg [7:0] out9047;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9047 = in0;
    end

    reg [7:0] out9048;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9048 = in0;
    end

    reg [7:0] out9049;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9049 = in0;
    end

    reg [7:0] out9050;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9050 = in0;
    end

    reg [7:0] out9051;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9051 = in0;
    end

    reg [7:0] out9052;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9052 = in0;
    end

    reg [7:0] out9053;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9053 = in0;
    end

    reg [7:0] out9054;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9054 = in0;
    end

    reg [7:0] out9055;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9055 = in0;
    end

    reg [7:0] out9056;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9056 = in0;
    end

    reg [7:0] out9057;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9057 = in0;
    end

    reg [7:0] out9058;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9058 = in0;
    end

    reg [7:0] out9059;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9059 = in0;
    end

    reg [7:0] out9060;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9060 = in0;
    end

    reg [7:0] out9061;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9061 = in0;
    end

    reg [7:0] out9062;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9062 = in0;
    end

    reg [7:0] out9063;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9063 = in0;
    end

    reg [7:0] out9064;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9064 = in0;
    end

    reg [7:0] out9065;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9065 = in0;
    end

    reg [7:0] out9066;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9066 = in0;
    end

    reg [7:0] out9067;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9067 = in0;
    end

    reg [7:0] out9068;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9068 = in0;
    end

    reg [7:0] out9069;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9069 = in0;
    end

    reg [7:0] out9070;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9070 = in0;
    end

    reg [7:0] out9071;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9071 = in0;
    end

    reg [7:0] out9072;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9072 = in0;
    end

    reg [7:0] out9073;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9073 = in0;
    end

    reg [7:0] out9074;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9074 = in0;
    end

    reg [7:0] out9075;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9075 = in0;
    end

    reg [7:0] out9076;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9076 = in0;
    end

    reg [7:0] out9077;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9077 = in0;
    end

    reg [7:0] out9078;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9078 = in0;
    end

    reg [7:0] out9079;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9079 = in0;
    end

    reg [7:0] out9080;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9080 = in0;
    end

    reg [7:0] out9081;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9081 = in0;
    end

    reg [7:0] out9082;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9082 = in0;
    end

    reg [7:0] out9083;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9083 = in0;
    end

    reg [7:0] out9084;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9084 = in0;
    end

    reg [7:0] out9085;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9085 = in0;
    end

    reg [7:0] out9086;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9086 = in0;
    end

    reg [7:0] out9087;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9087 = in0;
    end

    reg [7:0] out9088;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9088 = in0;
    end

    reg [7:0] out9089;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9089 = in0;
    end

    reg [7:0] out9090;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9090 = in0;
    end

    reg [7:0] out9091;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9091 = in0;
    end

    reg [7:0] out9092;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9092 = in0;
    end

    reg [7:0] out9093;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9093 = in0;
    end

    reg [7:0] out9094;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9094 = in0;
    end

    reg [7:0] out9095;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9095 = in0;
    end

    reg [7:0] out9096;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9096 = in0;
    end

    reg [7:0] out9097;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9097 = in0;
    end

    reg [7:0] out9098;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9098 = in0;
    end

    reg [7:0] out9099;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9099 = in0;
    end

    reg [7:0] out9100;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9100 = in0;
    end

    reg [7:0] out9101;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9101 = in0;
    end

    reg [7:0] out9102;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9102 = in0;
    end

    reg [7:0] out9103;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9103 = in0;
    end

    reg [7:0] out9104;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9104 = in0;
    end

    reg [7:0] out9105;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9105 = in0;
    end

    reg [7:0] out9106;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9106 = in0;
    end

    reg [7:0] out9107;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9107 = in0;
    end

    reg [7:0] out9108;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9108 = in0;
    end

    reg [7:0] out9109;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9109 = in0;
    end

    reg [7:0] out9110;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9110 = in0;
    end

    reg [7:0] out9111;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9111 = in0;
    end

    reg [7:0] out9112;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9112 = in0;
    end

    reg [7:0] out9113;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9113 = in0;
    end

    reg [7:0] out9114;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9114 = in0;
    end

    reg [7:0] out9115;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9115 = in0;
    end

    reg [7:0] out9116;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9116 = in0;
    end

    reg [7:0] out9117;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9117 = in0;
    end

    reg [7:0] out9118;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9118 = in0;
    end

    reg [7:0] out9119;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9119 = in0;
    end

    reg [7:0] out9120;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9120 = in0;
    end

    reg [7:0] out9121;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9121 = in0;
    end

    reg [7:0] out9122;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9122 = in0;
    end

    reg [7:0] out9123;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9123 = in0;
    end

    reg [7:0] out9124;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9124 = in0;
    end

    reg [7:0] out9125;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9125 = in0;
    end

    reg [7:0] out9126;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9126 = in0;
    end

    reg [7:0] out9127;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9127 = in0;
    end

    reg [7:0] out9128;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9128 = in0;
    end

    reg [7:0] out9129;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9129 = in0;
    end

    reg [7:0] out9130;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9130 = in0;
    end

    reg [7:0] out9131;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9131 = in0;
    end

    reg [7:0] out9132;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9132 = in0;
    end

    reg [7:0] out9133;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9133 = in0;
    end

    reg [7:0] out9134;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9134 = in0;
    end

    reg [7:0] out9135;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9135 = in0;
    end

    reg [7:0] out9136;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9136 = in0;
    end

    reg [7:0] out9137;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9137 = in0;
    end

    reg [7:0] out9138;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9138 = in0;
    end

    reg [7:0] out9139;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9139 = in0;
    end

    reg [7:0] out9140;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9140 = in0;
    end

    reg [7:0] out9141;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9141 = in0;
    end

    reg [7:0] out9142;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9142 = in0;
    end

    reg [7:0] out9143;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9143 = in0;
    end

    reg [7:0] out9144;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9144 = in0;
    end

    reg [7:0] out9145;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9145 = in0;
    end

    reg [7:0] out9146;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9146 = in0;
    end

    reg [7:0] out9147;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9147 = in0;
    end

    reg [7:0] out9148;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9148 = in0;
    end

    reg [7:0] out9149;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9149 = in0;
    end

    reg [7:0] out9150;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9150 = in0;
    end

    reg [7:0] out9151;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9151 = in0;
    end

    reg [7:0] out9152;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9152 = in0;
    end

    reg [7:0] out9153;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9153 = in0;
    end

    reg [7:0] out9154;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9154 = in0;
    end

    reg [7:0] out9155;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9155 = in0;
    end

    reg [7:0] out9156;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9156 = in0;
    end

    reg [7:0] out9157;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9157 = in0;
    end

    reg [7:0] out9158;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9158 = in0;
    end

    reg [7:0] out9159;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9159 = in0;
    end

    reg [7:0] out9160;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9160 = in0;
    end

    reg [7:0] out9161;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9161 = in0;
    end

    reg [7:0] out9162;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9162 = in0;
    end

    reg [7:0] out9163;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9163 = in0;
    end

    reg [7:0] out9164;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9164 = in0;
    end

    reg [7:0] out9165;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9165 = in0;
    end

    reg [7:0] out9166;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9166 = in0;
    end

    reg [7:0] out9167;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9167 = in0;
    end

    reg [7:0] out9168;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9168 = in0;
    end

    reg [7:0] out9169;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9169 = in0;
    end

    reg [7:0] out9170;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9170 = in0;
    end

    reg [7:0] out9171;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9171 = in0;
    end

    reg [7:0] out9172;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9172 = in0;
    end

    reg [7:0] out9173;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9173 = in0;
    end

    reg [7:0] out9174;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9174 = in0;
    end

    reg [7:0] out9175;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9175 = in0;
    end

    reg [7:0] out9176;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9176 = in0;
    end

    reg [7:0] out9177;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9177 = in0;
    end

    reg [7:0] out9178;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9178 = in0;
    end

    reg [7:0] out9179;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9179 = in0;
    end

    reg [7:0] out9180;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9180 = in0;
    end

    reg [7:0] out9181;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9181 = in0;
    end

    reg [7:0] out9182;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9182 = in0;
    end

    reg [7:0] out9183;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9183 = in0;
    end

    reg [7:0] out9184;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9184 = in0;
    end

    reg [7:0] out9185;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9185 = in0;
    end

    reg [7:0] out9186;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9186 = in0;
    end

    reg [7:0] out9187;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9187 = in0;
    end

    reg [7:0] out9188;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9188 = in0;
    end

    reg [7:0] out9189;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9189 = in0;
    end

    reg [7:0] out9190;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9190 = in0;
    end

    reg [7:0] out9191;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9191 = in0;
    end

    reg [7:0] out9192;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9192 = in0;
    end

    reg [7:0] out9193;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9193 = in0;
    end

    reg [7:0] out9194;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9194 = in0;
    end

    reg [7:0] out9195;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9195 = in0;
    end

    reg [7:0] out9196;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9196 = in0;
    end

    reg [7:0] out9197;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9197 = in0;
    end

    reg [7:0] out9198;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9198 = in0;
    end

    reg [7:0] out9199;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9199 = in0;
    end

    reg [7:0] out9200;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9200 = in0;
    end

    reg [7:0] out9201;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9201 = in0;
    end

    reg [7:0] out9202;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9202 = in0;
    end

    reg [7:0] out9203;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9203 = in0;
    end

    reg [7:0] out9204;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9204 = in0;
    end

    reg [7:0] out9205;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9205 = in0;
    end

    reg [7:0] out9206;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9206 = in0;
    end

    reg [7:0] out9207;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9207 = in0;
    end

    reg [7:0] out9208;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9208 = in0;
    end

    reg [7:0] out9209;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9209 = in0;
    end

    reg [7:0] out9210;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9210 = in0;
    end

    reg [7:0] out9211;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9211 = in0;
    end

    reg [7:0] out9212;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9212 = in0;
    end

    reg [7:0] out9213;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9213 = in0;
    end

    reg [7:0] out9214;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9214 = in0;
    end

    reg [7:0] out9215;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9215 = in0;
    end

    reg [7:0] out9216;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9216 = in0;
    end

    reg [7:0] out9217;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9217 = in0;
    end

    reg [7:0] out9218;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9218 = in0;
    end

    reg [7:0] out9219;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9219 = in0;
    end

    reg [7:0] out9220;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9220 = in0;
    end

    reg [7:0] out9221;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9221 = in0;
    end

    reg [7:0] out9222;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9222 = in0;
    end

    reg [7:0] out9223;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9223 = in0;
    end

    reg [7:0] out9224;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9224 = in0;
    end

    reg [7:0] out9225;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9225 = in0;
    end

    reg [7:0] out9226;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9226 = in0;
    end

    reg [7:0] out9227;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9227 = in0;
    end

    reg [7:0] out9228;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9228 = in0;
    end

    reg [7:0] out9229;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9229 = in0;
    end

    reg [7:0] out9230;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9230 = in0;
    end

    reg [7:0] out9231;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9231 = in0;
    end

    reg [7:0] out9232;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9232 = in0;
    end

    reg [7:0] out9233;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9233 = in0;
    end

    reg [7:0] out9234;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9234 = in0;
    end

    reg [7:0] out9235;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9235 = in0;
    end

    reg [7:0] out9236;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9236 = in0;
    end

    reg [7:0] out9237;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9237 = in0;
    end

    reg [7:0] out9238;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9238 = in0;
    end

    reg [7:0] out9239;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9239 = in0;
    end

    reg [7:0] out9240;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9240 = in0;
    end

    reg [7:0] out9241;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9241 = in0;
    end

    reg [7:0] out9242;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9242 = in0;
    end

    reg [7:0] out9243;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9243 = in0;
    end

    reg [7:0] out9244;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9244 = in0;
    end

    reg [7:0] out9245;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9245 = in0;
    end

    reg [7:0] out9246;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9246 = in0;
    end

    reg [7:0] out9247;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9247 = in0;
    end

    reg [7:0] out9248;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9248 = in0;
    end

    reg [7:0] out9249;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9249 = in0;
    end

    reg [7:0] out9250;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9250 = in0;
    end

    reg [7:0] out9251;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9251 = in0;
    end

    reg [7:0] out9252;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9252 = in0;
    end

    reg [7:0] out9253;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9253 = in0;
    end

    reg [7:0] out9254;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9254 = in0;
    end

    reg [7:0] out9255;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9255 = in0;
    end

    reg [7:0] out9256;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9256 = in0;
    end

    reg [7:0] out9257;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9257 = in0;
    end

    reg [7:0] out9258;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9258 = in0;
    end

    reg [7:0] out9259;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9259 = in0;
    end

    reg [7:0] out9260;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9260 = in0;
    end

    reg [7:0] out9261;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9261 = in0;
    end

    reg [7:0] out9262;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9262 = in0;
    end

    reg [7:0] out9263;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9263 = in0;
    end

    reg [7:0] out9264;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9264 = in0;
    end

    reg [7:0] out9265;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9265 = in0;
    end

    reg [7:0] out9266;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9266 = in0;
    end

    reg [7:0] out9267;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9267 = in0;
    end

    reg [7:0] out9268;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9268 = in0;
    end

    reg [7:0] out9269;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9269 = in0;
    end

    reg [7:0] out9270;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9270 = in0;
    end

    reg [7:0] out9271;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9271 = in0;
    end

    reg [7:0] out9272;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9272 = in0;
    end

    reg [7:0] out9273;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9273 = in0;
    end

    reg [7:0] out9274;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9274 = in0;
    end

    reg [7:0] out9275;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9275 = in0;
    end

    reg [7:0] out9276;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9276 = in0;
    end

    reg [7:0] out9277;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9277 = in0;
    end

    reg [7:0] out9278;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9278 = in0;
    end

    reg [7:0] out9279;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9279 = in0;
    end

    reg [7:0] out9280;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9280 = in0;
    end

    reg [7:0] out9281;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9281 = in0;
    end

    reg [7:0] out9282;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9282 = in0;
    end

    reg [7:0] out9283;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9283 = in0;
    end

    reg [7:0] out9284;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9284 = in0;
    end

    reg [7:0] out9285;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9285 = in0;
    end

    reg [7:0] out9286;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9286 = in0;
    end

    reg [7:0] out9287;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9287 = in0;
    end

    reg [7:0] out9288;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9288 = in0;
    end

    reg [7:0] out9289;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9289 = in0;
    end

    reg [7:0] out9290;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9290 = in0;
    end

    reg [7:0] out9291;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9291 = in0;
    end

    reg [7:0] out9292;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9292 = in0;
    end

    reg [7:0] out9293;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9293 = in0;
    end

    reg [7:0] out9294;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9294 = in0;
    end

    reg [7:0] out9295;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9295 = in0;
    end

    reg [7:0] out9296;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9296 = in0;
    end

    reg [7:0] out9297;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9297 = in0;
    end

    reg [7:0] out9298;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9298 = in0;
    end

    reg [7:0] out9299;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9299 = in0;
    end

    reg [7:0] out9300;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9300 = in0;
    end

    reg [7:0] out9301;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9301 = in0;
    end

    reg [7:0] out9302;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9302 = in0;
    end

    reg [7:0] out9303;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9303 = in0;
    end

    reg [7:0] out9304;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9304 = in0;
    end

    reg [7:0] out9305;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9305 = in0;
    end

    reg [7:0] out9306;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9306 = in0;
    end

    reg [7:0] out9307;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9307 = in0;
    end

    reg [7:0] out9308;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9308 = in0;
    end

    reg [7:0] out9309;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9309 = in0;
    end

    reg [7:0] out9310;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9310 = in0;
    end

    reg [7:0] out9311;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9311 = in0;
    end

    reg [7:0] out9312;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9312 = in0;
    end

    reg [7:0] out9313;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9313 = in0;
    end

    reg [7:0] out9314;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9314 = in0;
    end

    reg [7:0] out9315;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9315 = in0;
    end

    reg [7:0] out9316;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9316 = in0;
    end

    reg [7:0] out9317;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9317 = in0;
    end

    reg [7:0] out9318;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9318 = in0;
    end

    reg [7:0] out9319;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9319 = in0;
    end

    reg [7:0] out9320;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9320 = in0;
    end

    reg [7:0] out9321;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9321 = in0;
    end

    reg [7:0] out9322;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9322 = in0;
    end

    reg [7:0] out9323;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9323 = in0;
    end

    reg [7:0] out9324;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9324 = in0;
    end

    reg [7:0] out9325;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9325 = in0;
    end

    reg [7:0] out9326;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9326 = in0;
    end

    reg [7:0] out9327;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9327 = in0;
    end

    reg [7:0] out9328;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9328 = in0;
    end

    reg [7:0] out9329;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9329 = in0;
    end

    reg [7:0] out9330;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9330 = in0;
    end

    reg [7:0] out9331;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9331 = in0;
    end

    reg [7:0] out9332;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9332 = in0;
    end

    reg [7:0] out9333;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9333 = in0;
    end

    reg [7:0] out9334;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9334 = in0;
    end

    reg [7:0] out9335;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9335 = in0;
    end

    reg [7:0] out9336;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9336 = in0;
    end

    reg [7:0] out9337;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9337 = in0;
    end

    reg [7:0] out9338;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9338 = in0;
    end

    reg [7:0] out9339;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9339 = in0;
    end

    reg [7:0] out9340;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9340 = in0;
    end

    reg [7:0] out9341;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9341 = in0;
    end

    reg [7:0] out9342;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9342 = in0;
    end

    reg [7:0] out9343;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9343 = in0;
    end

    reg [7:0] out9344;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9344 = in0;
    end

    reg [7:0] out9345;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9345 = in0;
    end

    reg [7:0] out9346;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9346 = in0;
    end

    reg [7:0] out9347;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9347 = in0;
    end

    reg [7:0] out9348;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9348 = in0;
    end

    reg [7:0] out9349;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9349 = in0;
    end

    reg [7:0] out9350;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9350 = in0;
    end

    reg [7:0] out9351;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9351 = in0;
    end

    reg [7:0] out9352;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9352 = in0;
    end

    reg [7:0] out9353;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9353 = in0;
    end

    reg [7:0] out9354;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9354 = in0;
    end

    reg [7:0] out9355;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9355 = in0;
    end

    reg [7:0] out9356;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9356 = in0;
    end

    reg [7:0] out9357;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9357 = in0;
    end

    reg [7:0] out9358;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9358 = in0;
    end

    reg [7:0] out9359;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9359 = in0;
    end

    reg [7:0] out9360;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9360 = in0;
    end

    reg [7:0] out9361;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9361 = in0;
    end

    reg [7:0] out9362;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9362 = in0;
    end

    reg [7:0] out9363;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9363 = in0;
    end

    reg [7:0] out9364;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9364 = in0;
    end

    reg [7:0] out9365;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9365 = in0;
    end

    reg [7:0] out9366;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9366 = in0;
    end

    reg [7:0] out9367;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9367 = in0;
    end

    reg [7:0] out9368;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9368 = in0;
    end

    reg [7:0] out9369;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9369 = in0;
    end

    reg [7:0] out9370;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9370 = in0;
    end

    reg [7:0] out9371;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9371 = in0;
    end

    reg [7:0] out9372;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9372 = in0;
    end

    reg [7:0] out9373;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9373 = in0;
    end

    reg [7:0] out9374;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9374 = in0;
    end

    reg [7:0] out9375;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9375 = in0;
    end

    reg [7:0] out9376;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9376 = in0;
    end

    reg [7:0] out9377;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9377 = in0;
    end

    reg [7:0] out9378;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9378 = in0;
    end

    reg [7:0] out9379;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9379 = in0;
    end

    reg [7:0] out9380;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9380 = in0;
    end

    reg [7:0] out9381;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9381 = in0;
    end

    reg [7:0] out9382;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9382 = in0;
    end

    reg [7:0] out9383;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9383 = in0;
    end

    reg [7:0] out9384;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9384 = in0;
    end

    reg [7:0] out9385;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9385 = in0;
    end

    reg [7:0] out9386;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9386 = in0;
    end

    reg [7:0] out9387;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9387 = in0;
    end

    reg [7:0] out9388;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9388 = in0;
    end

    reg [7:0] out9389;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9389 = in0;
    end

    reg [7:0] out9390;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9390 = in0;
    end

    reg [7:0] out9391;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9391 = in0;
    end

    reg [7:0] out9392;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9392 = in0;
    end

    reg [7:0] out9393;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9393 = in0;
    end

    reg [7:0] out9394;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9394 = in0;
    end

    reg [7:0] out9395;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9395 = in0;
    end

    reg [7:0] out9396;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9396 = in0;
    end

    reg [7:0] out9397;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9397 = in0;
    end

    reg [7:0] out9398;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9398 = in0;
    end

    reg [7:0] out9399;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9399 = in0;
    end

    reg [7:0] out9400;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9400 = in0;
    end

    reg [7:0] out9401;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9401 = in0;
    end

    reg [7:0] out9402;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9402 = in0;
    end

    reg [7:0] out9403;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9403 = in0;
    end

    reg [7:0] out9404;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9404 = in0;
    end

    reg [7:0] out9405;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9405 = in0;
    end

    reg [7:0] out9406;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9406 = in0;
    end

    reg [7:0] out9407;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9407 = in0;
    end

    reg [7:0] out9408;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9408 = in0;
    end

    reg [7:0] out9409;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9409 = in0;
    end

    reg [7:0] out9410;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9410 = in0;
    end

    reg [7:0] out9411;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9411 = in0;
    end

    reg [7:0] out9412;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9412 = in0;
    end

    reg [7:0] out9413;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9413 = in0;
    end

    reg [7:0] out9414;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9414 = in0;
    end

    reg [7:0] out9415;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9415 = in0;
    end

    reg [7:0] out9416;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9416 = in0;
    end

    reg [7:0] out9417;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9417 = in0;
    end

    reg [7:0] out9418;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9418 = in0;
    end

    reg [7:0] out9419;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9419 = in0;
    end

    reg [7:0] out9420;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9420 = in0;
    end

    reg [7:0] out9421;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9421 = in0;
    end

    reg [7:0] out9422;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9422 = in0;
    end

    reg [7:0] out9423;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9423 = in0;
    end

    reg [7:0] out9424;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9424 = in0;
    end

    reg [7:0] out9425;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9425 = in0;
    end

    reg [7:0] out9426;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9426 = in0;
    end

    reg [7:0] out9427;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9427 = in0;
    end

    reg [7:0] out9428;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9428 = in0;
    end

    reg [7:0] out9429;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9429 = in0;
    end

    reg [7:0] out9430;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9430 = in0;
    end

    reg [7:0] out9431;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9431 = in0;
    end

    reg [7:0] out9432;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9432 = in0;
    end

    reg [7:0] out9433;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9433 = in0;
    end

    reg [7:0] out9434;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9434 = in0;
    end

    reg [7:0] out9435;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9435 = in0;
    end

    reg [7:0] out9436;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9436 = in0;
    end

    reg [7:0] out9437;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9437 = in0;
    end

    reg [7:0] out9438;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9438 = in0;
    end

    reg [7:0] out9439;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9439 = in0;
    end

    reg [7:0] out9440;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9440 = in0;
    end

    reg [7:0] out9441;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9441 = in0;
    end

    reg [7:0] out9442;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9442 = in0;
    end

    reg [7:0] out9443;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9443 = in0;
    end

    reg [7:0] out9444;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9444 = in0;
    end

    reg [7:0] out9445;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9445 = in0;
    end

    reg [7:0] out9446;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9446 = in0;
    end

    reg [7:0] out9447;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9447 = in0;
    end

    reg [7:0] out9448;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9448 = in0;
    end

    reg [7:0] out9449;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9449 = in0;
    end

    reg [7:0] out9450;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9450 = in0;
    end

    reg [7:0] out9451;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9451 = in0;
    end

    reg [7:0] out9452;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9452 = in0;
    end

    reg [7:0] out9453;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9453 = in0;
    end

    reg [7:0] out9454;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9454 = in0;
    end

    reg [7:0] out9455;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9455 = in0;
    end

    reg [7:0] out9456;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9456 = in0;
    end

    reg [7:0] out9457;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9457 = in0;
    end

    reg [7:0] out9458;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9458 = in0;
    end

    reg [7:0] out9459;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9459 = in0;
    end

    reg [7:0] out9460;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9460 = in0;
    end

    reg [7:0] out9461;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9461 = in0;
    end

    reg [7:0] out9462;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9462 = in0;
    end

    reg [7:0] out9463;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9463 = in0;
    end

    reg [7:0] out9464;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9464 = in0;
    end

    reg [7:0] out9465;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9465 = in0;
    end

    reg [7:0] out9466;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9466 = in0;
    end

    reg [7:0] out9467;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9467 = in0;
    end

    reg [7:0] out9468;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9468 = in0;
    end

    reg [7:0] out9469;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9469 = in0;
    end

    reg [7:0] out9470;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9470 = in0;
    end

    reg [7:0] out9471;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9471 = in0;
    end

    reg [7:0] out9472;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9472 = in0;
    end

    reg [7:0] out9473;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9473 = in0;
    end

    reg [7:0] out9474;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9474 = in0;
    end

    reg [7:0] out9475;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9475 = in0;
    end

    reg [7:0] out9476;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9476 = in0;
    end

    reg [7:0] out9477;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9477 = in0;
    end

    reg [7:0] out9478;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9478 = in0;
    end

    reg [7:0] out9479;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9479 = in0;
    end

    reg [7:0] out9480;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9480 = in0;
    end

    reg [7:0] out9481;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9481 = in0;
    end

    reg [7:0] out9482;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9482 = in0;
    end

    reg [7:0] out9483;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9483 = in0;
    end

    reg [7:0] out9484;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9484 = in0;
    end

    reg [7:0] out9485;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9485 = in0;
    end

    reg [7:0] out9486;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9486 = in0;
    end

    reg [7:0] out9487;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9487 = in0;
    end

    reg [7:0] out9488;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9488 = in0;
    end

    reg [7:0] out9489;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9489 = in0;
    end

    reg [7:0] out9490;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9490 = in0;
    end

    reg [7:0] out9491;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9491 = in0;
    end

    reg [7:0] out9492;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9492 = in0;
    end

    reg [7:0] out9493;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9493 = in0;
    end

    reg [7:0] out9494;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9494 = in0;
    end

    reg [7:0] out9495;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9495 = in0;
    end

    reg [7:0] out9496;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9496 = in0;
    end

    reg [7:0] out9497;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9497 = in0;
    end

    reg [7:0] out9498;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9498 = in0;
    end

    reg [7:0] out9499;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9499 = in0;
    end

    reg [7:0] out9500;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9500 = in0;
    end

    reg [7:0] out9501;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9501 = in0;
    end

    reg [7:0] out9502;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9502 = in0;
    end

    reg [7:0] out9503;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9503 = in0;
    end

    reg [7:0] out9504;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9504 = in0;
    end

    reg [7:0] out9505;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9505 = in0;
    end

    reg [7:0] out9506;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9506 = in0;
    end

    reg [7:0] out9507;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9507 = in0;
    end

    reg [7:0] out9508;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9508 = in0;
    end

    reg [7:0] out9509;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9509 = in0;
    end

    reg [7:0] out9510;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9510 = in0;
    end

    reg [7:0] out9511;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9511 = in0;
    end

    reg [7:0] out9512;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9512 = in0;
    end

    reg [7:0] out9513;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9513 = in0;
    end

    reg [7:0] out9514;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9514 = in0;
    end

    reg [7:0] out9515;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9515 = in0;
    end

    reg [7:0] out9516;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9516 = in0;
    end

    reg [7:0] out9517;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9517 = in0;
    end

    reg [7:0] out9518;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9518 = in0;
    end

    reg [7:0] out9519;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9519 = in0;
    end

    reg [7:0] out9520;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9520 = in0;
    end

    reg [7:0] out9521;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9521 = in0;
    end

    reg [7:0] out9522;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9522 = in0;
    end

    reg [7:0] out9523;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9523 = in0;
    end

    reg [7:0] out9524;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9524 = in0;
    end

    reg [7:0] out9525;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9525 = in0;
    end

    reg [7:0] out9526;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9526 = in0;
    end

    reg [7:0] out9527;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9527 = in0;
    end

    reg [7:0] out9528;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9528 = in0;
    end

    reg [7:0] out9529;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9529 = in0;
    end

    reg [7:0] out9530;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9530 = in0;
    end

    reg [7:0] out9531;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9531 = in0;
    end

    reg [7:0] out9532;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9532 = in0;
    end

    reg [7:0] out9533;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9533 = in0;
    end

    reg [7:0] out9534;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9534 = in0;
    end

    reg [7:0] out9535;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9535 = in0;
    end

    reg [7:0] out9536;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9536 = in0;
    end

    reg [7:0] out9537;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9537 = in0;
    end

    reg [7:0] out9538;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9538 = in0;
    end

    reg [7:0] out9539;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9539 = in0;
    end

    reg [7:0] out9540;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9540 = in0;
    end

    reg [7:0] out9541;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9541 = in0;
    end

    reg [7:0] out9542;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9542 = in0;
    end

    reg [7:0] out9543;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9543 = in0;
    end

    reg [7:0] out9544;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9544 = in0;
    end

    reg [7:0] out9545;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9545 = in0;
    end

    reg [7:0] out9546;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9546 = in0;
    end

    reg [7:0] out9547;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9547 = in0;
    end

    reg [7:0] out9548;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9548 = in0;
    end

    reg [7:0] out9549;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9549 = in0;
    end

    reg [7:0] out9550;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9550 = in0;
    end

    reg [7:0] out9551;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9551 = in0;
    end

    reg [7:0] out9552;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9552 = in0;
    end

    reg [7:0] out9553;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9553 = in0;
    end

    reg [7:0] out9554;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9554 = in0;
    end

    reg [7:0] out9555;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9555 = in0;
    end

    reg [7:0] out9556;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9556 = in0;
    end

    reg [7:0] out9557;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9557 = in0;
    end

    reg [7:0] out9558;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9558 = in0;
    end

    reg [7:0] out9559;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9559 = in0;
    end

    reg [7:0] out9560;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9560 = in0;
    end

    reg [7:0] out9561;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9561 = in0;
    end

    reg [7:0] out9562;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9562 = in0;
    end

    reg [7:0] out9563;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9563 = in0;
    end

    reg [7:0] out9564;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9564 = in0;
    end

    reg [7:0] out9565;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9565 = in0;
    end

    reg [7:0] out9566;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9566 = in0;
    end

    reg [7:0] out9567;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9567 = in0;
    end

    reg [7:0] out9568;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9568 = in0;
    end

    reg [7:0] out9569;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9569 = in0;
    end

    reg [7:0] out9570;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9570 = in0;
    end

    reg [7:0] out9571;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9571 = in0;
    end

    reg [7:0] out9572;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9572 = in0;
    end

    reg [7:0] out9573;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9573 = in0;
    end

    reg [7:0] out9574;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9574 = in0;
    end

    reg [7:0] out9575;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9575 = in0;
    end

    reg [7:0] out9576;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9576 = in0;
    end

    reg [7:0] out9577;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9577 = in0;
    end

    reg [7:0] out9578;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9578 = in0;
    end

    reg [7:0] out9579;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9579 = in0;
    end

    reg [7:0] out9580;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9580 = in0;
    end

    reg [7:0] out9581;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9581 = in0;
    end

    reg [7:0] out9582;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9582 = in0;
    end

    reg [7:0] out9583;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9583 = in0;
    end

    reg [7:0] out9584;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9584 = in0;
    end

    reg [7:0] out9585;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9585 = in0;
    end

    reg [7:0] out9586;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9586 = in0;
    end

    reg [7:0] out9587;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9587 = in0;
    end

    reg [7:0] out9588;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9588 = in0;
    end

    reg [7:0] out9589;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9589 = in0;
    end

    reg [7:0] out9590;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9590 = in0;
    end

    reg [7:0] out9591;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9591 = in0;
    end

    reg [7:0] out9592;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9592 = in0;
    end

    reg [7:0] out9593;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9593 = in0;
    end

    reg [7:0] out9594;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9594 = in0;
    end

    reg [7:0] out9595;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9595 = in0;
    end

    reg [7:0] out9596;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9596 = in0;
    end

    reg [7:0] out9597;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9597 = in0;
    end

    reg [7:0] out9598;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9598 = in0;
    end

    reg [7:0] out9599;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9599 = in0;
    end

    reg [7:0] out9600;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9600 = in0;
    end

    reg [7:0] out9601;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9601 = in0;
    end

    reg [7:0] out9602;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9602 = in0;
    end

    reg [7:0] out9603;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9603 = in0;
    end

    reg [7:0] out9604;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9604 = in0;
    end

    reg [7:0] out9605;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9605 = in0;
    end

    reg [7:0] out9606;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9606 = in0;
    end

    reg [7:0] out9607;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9607 = in0;
    end

    reg [7:0] out9608;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9608 = in0;
    end

    reg [7:0] out9609;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9609 = in0;
    end

    reg [7:0] out9610;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9610 = in0;
    end

    reg [7:0] out9611;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9611 = in0;
    end

    reg [7:0] out9612;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9612 = in0;
    end

    reg [7:0] out9613;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9613 = in0;
    end

    reg [7:0] out9614;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9614 = in0;
    end

    reg [7:0] out9615;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9615 = in0;
    end

    reg [7:0] out9616;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9616 = in0;
    end

    reg [7:0] out9617;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9617 = in0;
    end

    reg [7:0] out9618;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9618 = in0;
    end

    reg [7:0] out9619;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9619 = in0;
    end

    reg [7:0] out9620;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9620 = in0;
    end

    reg [7:0] out9621;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9621 = in0;
    end

    reg [7:0] out9622;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9622 = in0;
    end

    reg [7:0] out9623;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9623 = in0;
    end

    reg [7:0] out9624;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9624 = in0;
    end

    reg [7:0] out9625;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9625 = in0;
    end

    reg [7:0] out9626;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9626 = in0;
    end

    reg [7:0] out9627;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9627 = in0;
    end

    reg [7:0] out9628;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9628 = in0;
    end

    reg [7:0] out9629;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9629 = in0;
    end

    reg [7:0] out9630;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9630 = in0;
    end

    reg [7:0] out9631;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9631 = in0;
    end

    reg [7:0] out9632;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9632 = in0;
    end

    reg [7:0] out9633;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9633 = in0;
    end

    reg [7:0] out9634;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9634 = in0;
    end

    reg [7:0] out9635;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9635 = in0;
    end

    reg [7:0] out9636;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9636 = in0;
    end

    reg [7:0] out9637;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9637 = in0;
    end

    reg [7:0] out9638;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9638 = in0;
    end

    reg [7:0] out9639;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9639 = in0;
    end

    reg [7:0] out9640;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9640 = in0;
    end

    reg [7:0] out9641;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9641 = in0;
    end

    reg [7:0] out9642;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9642 = in0;
    end

    reg [7:0] out9643;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9643 = in0;
    end

    reg [7:0] out9644;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9644 = in0;
    end

    reg [7:0] out9645;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9645 = in0;
    end

    reg [7:0] out9646;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9646 = in0;
    end

    reg [7:0] out9647;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9647 = in0;
    end

    reg [7:0] out9648;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9648 = in0;
    end

    reg [7:0] out9649;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9649 = in0;
    end

    reg [7:0] out9650;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9650 = in0;
    end

    reg [7:0] out9651;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9651 = in0;
    end

    reg [7:0] out9652;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9652 = in0;
    end

    reg [7:0] out9653;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9653 = in0;
    end

    reg [7:0] out9654;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9654 = in0;
    end

    reg [7:0] out9655;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9655 = in0;
    end

    reg [7:0] out9656;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9656 = in0;
    end

    reg [7:0] out9657;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9657 = in0;
    end

    reg [7:0] out9658;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9658 = in0;
    end

    reg [7:0] out9659;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9659 = in0;
    end

    reg [7:0] out9660;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9660 = in0;
    end

    reg [7:0] out9661;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9661 = in0;
    end

    reg [7:0] out9662;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9662 = in0;
    end

    reg [7:0] out9663;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9663 = in0;
    end

    reg [7:0] out9664;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9664 = in0;
    end

    reg [7:0] out9665;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9665 = in0;
    end

    reg [7:0] out9666;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9666 = in0;
    end

    reg [7:0] out9667;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9667 = in0;
    end

    reg [7:0] out9668;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9668 = in0;
    end

    reg [7:0] out9669;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9669 = in0;
    end

    reg [7:0] out9670;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9670 = in0;
    end

    reg [7:0] out9671;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9671 = in0;
    end

    reg [7:0] out9672;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9672 = in0;
    end

    reg [7:0] out9673;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9673 = in0;
    end

    reg [7:0] out9674;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9674 = in0;
    end

    reg [7:0] out9675;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9675 = in0;
    end

    reg [7:0] out9676;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9676 = in0;
    end

    reg [7:0] out9677;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9677 = in0;
    end

    reg [7:0] out9678;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9678 = in0;
    end

    reg [7:0] out9679;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9679 = in0;
    end

    reg [7:0] out9680;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9680 = in0;
    end

    reg [7:0] out9681;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9681 = in0;
    end

    reg [7:0] out9682;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9682 = in0;
    end

    reg [7:0] out9683;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9683 = in0;
    end

    reg [7:0] out9684;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9684 = in0;
    end

    reg [7:0] out9685;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9685 = in0;
    end

    reg [7:0] out9686;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9686 = in0;
    end

    reg [7:0] out9687;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9687 = in0;
    end

    reg [7:0] out9688;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9688 = in0;
    end

    reg [7:0] out9689;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9689 = in0;
    end

    reg [7:0] out9690;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9690 = in0;
    end

    reg [7:0] out9691;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9691 = in0;
    end

    reg [7:0] out9692;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9692 = in0;
    end

    reg [7:0] out9693;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9693 = in0;
    end

    reg [7:0] out9694;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9694 = in0;
    end

    reg [7:0] out9695;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9695 = in0;
    end

    reg [7:0] out9696;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9696 = in0;
    end

    reg [7:0] out9697;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9697 = in0;
    end

    reg [7:0] out9698;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9698 = in0;
    end

    reg [7:0] out9699;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9699 = in0;
    end

    reg [7:0] out9700;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9700 = in0;
    end

    reg [7:0] out9701;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9701 = in0;
    end

    reg [7:0] out9702;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9702 = in0;
    end

    reg [7:0] out9703;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9703 = in0;
    end

    reg [7:0] out9704;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9704 = in0;
    end

    reg [7:0] out9705;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9705 = in0;
    end

    reg [7:0] out9706;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9706 = in0;
    end

    reg [7:0] out9707;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9707 = in0;
    end

    reg [7:0] out9708;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9708 = in0;
    end

    reg [7:0] out9709;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9709 = in0;
    end

    reg [7:0] out9710;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9710 = in0;
    end

    reg [7:0] out9711;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9711 = in0;
    end

    reg [7:0] out9712;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9712 = in0;
    end

    reg [7:0] out9713;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9713 = in0;
    end

    reg [7:0] out9714;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9714 = in0;
    end

    reg [7:0] out9715;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9715 = in0;
    end

    reg [7:0] out9716;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9716 = in0;
    end

    reg [7:0] out9717;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9717 = in0;
    end

    reg [7:0] out9718;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9718 = in0;
    end

    reg [7:0] out9719;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9719 = in0;
    end

    reg [7:0] out9720;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9720 = in0;
    end

    reg [7:0] out9721;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9721 = in0;
    end

    reg [7:0] out9722;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9722 = in0;
    end

    reg [7:0] out9723;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9723 = in0;
    end

    reg [7:0] out9724;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9724 = in0;
    end

    reg [7:0] out9725;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9725 = in0;
    end

    reg [7:0] out9726;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9726 = in0;
    end

    reg [7:0] out9727;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9727 = in0;
    end

    reg [7:0] out9728;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9728 = in0;
    end

    reg [7:0] out9729;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9729 = in0;
    end

    reg [7:0] out9730;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9730 = in0;
    end

    reg [7:0] out9731;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9731 = in0;
    end

    reg [7:0] out9732;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9732 = in0;
    end

    reg [7:0] out9733;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9733 = in0;
    end

    reg [7:0] out9734;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9734 = in0;
    end

    reg [7:0] out9735;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9735 = in0;
    end

    reg [7:0] out9736;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9736 = in0;
    end

    reg [7:0] out9737;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9737 = in0;
    end

    reg [7:0] out9738;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9738 = in0;
    end

    reg [7:0] out9739;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9739 = in0;
    end

    reg [7:0] out9740;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9740 = in0;
    end

    reg [7:0] out9741;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9741 = in0;
    end

    reg [7:0] out9742;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9742 = in0;
    end

    reg [7:0] out9743;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9743 = in0;
    end

    reg [7:0] out9744;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9744 = in0;
    end

    reg [7:0] out9745;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9745 = in0;
    end

    reg [7:0] out9746;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9746 = in0;
    end

    reg [7:0] out9747;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9747 = in0;
    end

    reg [7:0] out9748;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9748 = in0;
    end

    reg [7:0] out9749;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9749 = in0;
    end

    reg [7:0] out9750;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9750 = in0;
    end

    reg [7:0] out9751;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9751 = in0;
    end

    reg [7:0] out9752;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9752 = in0;
    end

    reg [7:0] out9753;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9753 = in0;
    end

    reg [7:0] out9754;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9754 = in0;
    end

    reg [7:0] out9755;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9755 = in0;
    end

    reg [7:0] out9756;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9756 = in0;
    end

    reg [7:0] out9757;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9757 = in0;
    end

    reg [7:0] out9758;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9758 = in0;
    end

    reg [7:0] out9759;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9759 = in0;
    end

    reg [7:0] out9760;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9760 = in0;
    end

    reg [7:0] out9761;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9761 = in0;
    end

    reg [7:0] out9762;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9762 = in0;
    end

    reg [7:0] out9763;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9763 = in0;
    end

    reg [7:0] out9764;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9764 = in0;
    end

    reg [7:0] out9765;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9765 = in0;
    end

    reg [7:0] out9766;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9766 = in0;
    end

    reg [7:0] out9767;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9767 = in0;
    end

    reg [7:0] out9768;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9768 = in0;
    end

    reg [7:0] out9769;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9769 = in0;
    end

    reg [7:0] out9770;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9770 = in0;
    end

    reg [7:0] out9771;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9771 = in0;
    end

    reg [7:0] out9772;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9772 = in0;
    end

    reg [7:0] out9773;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9773 = in0;
    end

    reg [7:0] out9774;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9774 = in0;
    end

    reg [7:0] out9775;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9775 = in0;
    end

    reg [7:0] out9776;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9776 = in0;
    end

    reg [7:0] out9777;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9777 = in0;
    end

    reg [7:0] out9778;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9778 = in0;
    end

    reg [7:0] out9779;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9779 = in0;
    end

    reg [7:0] out9780;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9780 = in0;
    end

    reg [7:0] out9781;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9781 = in0;
    end

    reg [7:0] out9782;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9782 = in0;
    end

    reg [7:0] out9783;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9783 = in0;
    end

    reg [7:0] out9784;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9784 = in0;
    end

    reg [7:0] out9785;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9785 = in0;
    end

    reg [7:0] out9786;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9786 = in0;
    end

    reg [7:0] out9787;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9787 = in0;
    end

    reg [7:0] out9788;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9788 = in0;
    end

    reg [7:0] out9789;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9789 = in0;
    end

    reg [7:0] out9790;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9790 = in0;
    end

    reg [7:0] out9791;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9791 = in0;
    end

    reg [7:0] out9792;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9792 = in0;
    end

    reg [7:0] out9793;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9793 = in0;
    end

    reg [7:0] out9794;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9794 = in0;
    end

    reg [7:0] out9795;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9795 = in0;
    end

    reg [7:0] out9796;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9796 = in0;
    end

    reg [7:0] out9797;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9797 = in0;
    end

    reg [7:0] out9798;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9798 = in0;
    end

    reg [7:0] out9799;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9799 = in0;
    end

    reg [7:0] out9800;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9800 = in0;
    end

    reg [7:0] out9801;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9801 = in0;
    end

    reg [7:0] out9802;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9802 = in0;
    end

    reg [7:0] out9803;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9803 = in0;
    end

    reg [7:0] out9804;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9804 = in0;
    end

    reg [7:0] out9805;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9805 = in0;
    end

    reg [7:0] out9806;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9806 = in0;
    end

    reg [7:0] out9807;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9807 = in0;
    end

    reg [7:0] out9808;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9808 = in0;
    end

    reg [7:0] out9809;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9809 = in0;
    end

    reg [7:0] out9810;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9810 = in0;
    end

    reg [7:0] out9811;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9811 = in0;
    end

    reg [7:0] out9812;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9812 = in0;
    end

    reg [7:0] out9813;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9813 = in0;
    end

    reg [7:0] out9814;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9814 = in0;
    end

    reg [7:0] out9815;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9815 = in0;
    end

    reg [7:0] out9816;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9816 = in0;
    end

    reg [7:0] out9817;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9817 = in0;
    end

    reg [7:0] out9818;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9818 = in0;
    end

    reg [7:0] out9819;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9819 = in0;
    end

    reg [7:0] out9820;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9820 = in0;
    end

    reg [7:0] out9821;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9821 = in0;
    end

    reg [7:0] out9822;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9822 = in0;
    end

    reg [7:0] out9823;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9823 = in0;
    end

    reg [7:0] out9824;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9824 = in0;
    end

    reg [7:0] out9825;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9825 = in0;
    end

    reg [7:0] out9826;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9826 = in0;
    end

    reg [7:0] out9827;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9827 = in0;
    end

    reg [7:0] out9828;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9828 = in0;
    end

    reg [7:0] out9829;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9829 = in0;
    end

    reg [7:0] out9830;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9830 = in0;
    end

    reg [7:0] out9831;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9831 = in0;
    end

    reg [7:0] out9832;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9832 = in0;
    end

    reg [7:0] out9833;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9833 = in0;
    end

    reg [7:0] out9834;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9834 = in0;
    end

    reg [7:0] out9835;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9835 = in0;
    end

    reg [7:0] out9836;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9836 = in0;
    end

    reg [7:0] out9837;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9837 = in0;
    end

    reg [7:0] out9838;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9838 = in0;
    end

    reg [7:0] out9839;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9839 = in0;
    end

    reg [7:0] out9840;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9840 = in0;
    end

    reg [7:0] out9841;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9841 = in0;
    end

    reg [7:0] out9842;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9842 = in0;
    end

    reg [7:0] out9843;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9843 = in0;
    end

    reg [7:0] out9844;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9844 = in0;
    end

    reg [7:0] out9845;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9845 = in0;
    end

    reg [7:0] out9846;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9846 = in0;
    end

    reg [7:0] out9847;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9847 = in0;
    end

    reg [7:0] out9848;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9848 = in0;
    end

    reg [7:0] out9849;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9849 = in0;
    end

    reg [7:0] out9850;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9850 = in0;
    end

    reg [7:0] out9851;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9851 = in0;
    end

    reg [7:0] out9852;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9852 = in0;
    end

    reg [7:0] out9853;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9853 = in0;
    end

    reg [7:0] out9854;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9854 = in0;
    end

    reg [7:0] out9855;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9855 = in0;
    end

    reg [7:0] out9856;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9856 = in0;
    end

    reg [7:0] out9857;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9857 = in0;
    end

    reg [7:0] out9858;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9858 = in0;
    end

    reg [7:0] out9859;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9859 = in0;
    end

    reg [7:0] out9860;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9860 = in0;
    end

    reg [7:0] out9861;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9861 = in0;
    end

    reg [7:0] out9862;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9862 = in0;
    end

    reg [7:0] out9863;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9863 = in0;
    end

    reg [7:0] out9864;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9864 = in0;
    end

    reg [7:0] out9865;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9865 = in0;
    end

    reg [7:0] out9866;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9866 = in0;
    end

    reg [7:0] out9867;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9867 = in0;
    end

    reg [7:0] out9868;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9868 = in0;
    end

    reg [7:0] out9869;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9869 = in0;
    end

    reg [7:0] out9870;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9870 = in0;
    end

    reg [7:0] out9871;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9871 = in0;
    end

    reg [7:0] out9872;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9872 = in0;
    end

    reg [7:0] out9873;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9873 = in0;
    end

    reg [7:0] out9874;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9874 = in0;
    end

    reg [7:0] out9875;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9875 = in0;
    end

    reg [7:0] out9876;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9876 = in0;
    end

    reg [7:0] out9877;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9877 = in0;
    end

    reg [7:0] out9878;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9878 = in0;
    end

    reg [7:0] out9879;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9879 = in0;
    end

    reg [7:0] out9880;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9880 = in0;
    end

    reg [7:0] out9881;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9881 = in0;
    end

    reg [7:0] out9882;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9882 = in0;
    end

    reg [7:0] out9883;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9883 = in0;
    end

    reg [7:0] out9884;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9884 = in0;
    end

    reg [7:0] out9885;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9885 = in0;
    end

    reg [7:0] out9886;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9886 = in0;
    end

    reg [7:0] out9887;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9887 = in0;
    end

    reg [7:0] out9888;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9888 = in0;
    end

    reg [7:0] out9889;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9889 = in0;
    end

    reg [7:0] out9890;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9890 = in0;
    end

    reg [7:0] out9891;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9891 = in0;
    end

    reg [7:0] out9892;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9892 = in0;
    end

    reg [7:0] out9893;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9893 = in0;
    end

    reg [7:0] out9894;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9894 = in0;
    end

    reg [7:0] out9895;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9895 = in0;
    end

    reg [7:0] out9896;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9896 = in0;
    end

    reg [7:0] out9897;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9897 = in0;
    end

    reg [7:0] out9898;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9898 = in0;
    end

    reg [7:0] out9899;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9899 = in0;
    end

    reg [7:0] out9900;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9900 = in0;
    end

    reg [7:0] out9901;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9901 = in0;
    end

    reg [7:0] out9902;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9902 = in0;
    end

    reg [7:0] out9903;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9903 = in0;
    end

    reg [7:0] out9904;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9904 = in0;
    end

    reg [7:0] out9905;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9905 = in0;
    end

    reg [7:0] out9906;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9906 = in0;
    end

    reg [7:0] out9907;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9907 = in0;
    end

    reg [7:0] out9908;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9908 = in0;
    end

    reg [7:0] out9909;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9909 = in0;
    end

    reg [7:0] out9910;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9910 = in0;
    end

    reg [7:0] out9911;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9911 = in0;
    end

    reg [7:0] out9912;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9912 = in0;
    end

    reg [7:0] out9913;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9913 = in0;
    end

    reg [7:0] out9914;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9914 = in0;
    end

    reg [7:0] out9915;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9915 = in0;
    end

    reg [7:0] out9916;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9916 = in0;
    end

    reg [7:0] out9917;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9917 = in0;
    end

    reg [7:0] out9918;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9918 = in0;
    end

    reg [7:0] out9919;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9919 = in0;
    end

    reg [7:0] out9920;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9920 = in0;
    end

    reg [7:0] out9921;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9921 = in0;
    end

    reg [7:0] out9922;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9922 = in0;
    end

    reg [7:0] out9923;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9923 = in0;
    end

    reg [7:0] out9924;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9924 = in0;
    end

    reg [7:0] out9925;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9925 = in0;
    end

    reg [7:0] out9926;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9926 = in0;
    end

    reg [7:0] out9927;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9927 = in0;
    end

    reg [7:0] out9928;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9928 = in0;
    end

    reg [7:0] out9929;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9929 = in0;
    end

    reg [7:0] out9930;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9930 = in0;
    end

    reg [7:0] out9931;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9931 = in0;
    end

    reg [7:0] out9932;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9932 = in0;
    end

    reg [7:0] out9933;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9933 = in0;
    end

    reg [7:0] out9934;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9934 = in0;
    end

    reg [7:0] out9935;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9935 = in0;
    end

    reg [7:0] out9936;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9936 = in0;
    end

    reg [7:0] out9937;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9937 = in0;
    end

    reg [7:0] out9938;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9938 = in0;
    end

    reg [7:0] out9939;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9939 = in0;
    end

    reg [7:0] out9940;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9940 = in0;
    end

    reg [7:0] out9941;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9941 = in0;
    end

    reg [7:0] out9942;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9942 = in0;
    end

    reg [7:0] out9943;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9943 = in0;
    end

    reg [7:0] out9944;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9944 = in0;
    end

    reg [7:0] out9945;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9945 = in0;
    end

    reg [7:0] out9946;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9946 = in0;
    end

    reg [7:0] out9947;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9947 = in0;
    end

    reg [7:0] out9948;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9948 = in0;
    end

    reg [7:0] out9949;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9949 = in0;
    end

    reg [7:0] out9950;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9950 = in0;
    end

    reg [7:0] out9951;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9951 = in0;
    end

    reg [7:0] out9952;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9952 = in0;
    end

    reg [7:0] out9953;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9953 = in0;
    end

    reg [7:0] out9954;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9954 = in0;
    end

    reg [7:0] out9955;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9955 = in0;
    end

    reg [7:0] out9956;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9956 = in0;
    end

    reg [7:0] out9957;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9957 = in0;
    end

    reg [7:0] out9958;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9958 = in0;
    end

    reg [7:0] out9959;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9959 = in0;
    end

    reg [7:0] out9960;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9960 = in0;
    end

    reg [7:0] out9961;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9961 = in0;
    end

    reg [7:0] out9962;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9962 = in0;
    end

    reg [7:0] out9963;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9963 = in0;
    end

    reg [7:0] out9964;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9964 = in0;
    end

    reg [7:0] out9965;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9965 = in0;
    end

    reg [7:0] out9966;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9966 = in0;
    end

    reg [7:0] out9967;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9967 = in0;
    end

    reg [7:0] out9968;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9968 = in0;
    end

    reg [7:0] out9969;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9969 = in0;
    end

    reg [7:0] out9970;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9970 = in0;
    end

    reg [7:0] out9971;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9971 = in0;
    end

    reg [7:0] out9972;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9972 = in0;
    end

    reg [7:0] out9973;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9973 = in0;
    end

    reg [7:0] out9974;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9974 = in0;
    end

    reg [7:0] out9975;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9975 = in0;
    end

    reg [7:0] out9976;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9976 = in0;
    end

    reg [7:0] out9977;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9977 = in0;
    end

    reg [7:0] out9978;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9978 = in0;
    end

    reg [7:0] out9979;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9979 = in0;
    end

    reg [7:0] out9980;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9980 = in0;
    end

    reg [7:0] out9981;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9981 = in0;
    end

    reg [7:0] out9982;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9982 = in0;
    end

    reg [7:0] out9983;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9983 = in0;
    end

    reg [7:0] out9984;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9984 = in0;
    end

    reg [7:0] out9985;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9985 = in0;
    end

    reg [7:0] out9986;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9986 = in0;
    end

    reg [7:0] out9987;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9987 = in0;
    end

    reg [7:0] out9988;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9988 = in0;
    end

    reg [7:0] out9989;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9989 = in0;
    end

    reg [7:0] out9990;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9990 = in0;
    end

    reg [7:0] out9991;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9991 = in0;
    end

    reg [7:0] out9992;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9992 = in0;
    end

    reg [7:0] out9993;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9993 = in0;
    end

    reg [7:0] out9994;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9994 = in0;
    end

    reg [7:0] out9995;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9995 = in0;
    end

    reg [7:0] out9996;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9996 = in0;
    end

    reg [7:0] out9997;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9997 = in0;
    end

    reg [7:0] out9998;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9998 = in0;
    end

    reg [7:0] out9999;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out9999 = in0;
    end

    reg [7:0] out10000;

    always @(in0)
    for(i = 0;i<8;i++) begin
        out10000 = in0;
    end

    initial begin
        out1 = 0;
    end

    initial begin
        out2 = 0;
    end

    initial begin
        out3 = 0;
    end

    initial begin
        out4 = 0;
    end

    initial begin
        out5 = 0;
    end

    initial begin
        out6 = 0;
    end

    initial begin
        out7 = 0;
    end

    initial begin
        out8 = 0;
    end

    initial begin
        out9 = 0;
    end

    initial begin
        out10 = 0;
    end
endmodule
